library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"91",X"50",X"2F",X"4D",X"DE",X"81",X"A0",X"88",X"82",X"90",X"28",X"EB",X"FC",X"8B",X"88",X"A0",
		X"B2",X"48",X"18",X"0F",X"00",X"08",X"2F",X"5E",X"07",X"08",X"A8",X"2F",X"77",X"61",X"CD",X"BB",
		X"A0",X"C9",X"69",X"16",X"5F",X"D7",X"41",X"69",X"A0",X"88",X"A0",X"88",X"A0",X"88",X"A0",X"88",
		X"28",X"88",X"28",X"88",X"28",X"88",X"28",X"88",X"A8",X"71",X"DD",X"ED",X"D5",X"ED",X"A2",X"88",
		X"28",X"CD",X"B2",X"8A",X"28",X"DD",X"27",X"92",X"D0",X"18",X"92",X"C8",X"B8",X"12",X"80",X"28",
		X"07",X"08",X"2C",X"1D",X"32",X"80",X"88",X"1A",X"21",X"28",X"07",X"08",X"2C",X"1D",X"32",X"81",
		X"28",X"12",X"5F",X"0F",X"07",X"EA",X"17",X"89",X"A2",X"82",X"28",X"83",X"82",X"82",X"28",X"6D",
		X"94",X"92",X"CD",X"02",X"2A",X"65",X"CD",X"8A",X"CD",X"F7",X"2A",X"65",X"12",X"8B",X"CD",X"22",
		X"A3",X"81",X"73",X"2C",X"94",X"16",X"15",X"1E",X"90",X"9C",X"96",X"88",X"83",X"94",X"B6",X"B3",
		X"96",X"98",X"AB",X"9E",X"28",X"8B",X"34",X"3E",X"30",X"8C",X"36",X"88",X"23",X"9C",X"B6",X"88",
		X"7D",X"81",X"C0",X"2C",X"6D",X"39",X"32",X"16",X"A1",X"7D",X"81",X"D0",X"2C",X"6D",X"39",X"BA",
		X"B6",X"8B",X"DD",X"89",X"18",X"2C",X"CD",X"39",X"BA",X"1E",X"2A",X"75",X"21",X"08",X"8C",X"65",
		X"39",X"BA",X"B6",X"8C",X"7D",X"81",X"88",X"2C",X"6D",X"39",X"32",X"81",X"80",X"2F",X"B2",X"34",
		X"8C",X"AF",X"A0",X"8B",X"21",X"A0",X"8F",X"91",X"2E",X"2F",X"29",X"8D",X"28",X"6D",X"10",X"5E",
		X"92",X"99",X"2F",X"81",X"90",X"2F",X"B2",X"35",X"2C",X"8F",X"A0",X"8B",X"81",X"B0",X"2F",X"B1",
		X"AB",X"2F",X"29",X"8D",X"28",X"6D",X"10",X"5E",X"32",X"9A",X"8F",X"89",X"97",X"2C",X"CB",X"C6",
		X"80",X"05",X"63",X"0E",X"89",X"08",X"2F",X"39",X"B0",X"38",X"09",X"18",X"A0",X"C5",X"B8",X"B2",
		X"38",X"8F",X"CB",X"F7",X"A0",X"08",X"46",X"07",X"32",X"10",X"8F",X"32",X"2D",X"90",X"B2",X"11",
		X"2F",X"CB",X"D7",X"A0",X"20",X"46",X"A7",X"32",X"B1",X"27",X"9A",X"02",X"B8",X"B2",X"B2",X"27",
		X"CB",X"F7",X"A0",X"08",X"46",X"07",X"32",X"12",X"8F",X"32",X"AF",X"90",X"CD",X"94",X"29",X"51",
		X"9A",X"0A",X"28",X"41",X"8A",X"08",X"28",X"D5",X"E9",X"DD",X"E9",X"D9",X"65",X"53",X"A1",X"CD",
		X"F1",X"01",X"B6",X"01",X"32",X"40",X"18",X"A8",X"D3",X"C5",X"ED",X"B2",X"B9",X"88",X"07",X"48",
		X"92",X"00",X"28",X"07",X"60",X"B6",X"A1",X"32",X"31",X"20",X"99",X"F8",X"2F",X"21",X"B8",X"0C",
		X"45",X"B6",X"29",X"32",X"68",X"90",X"D3",X"C5",X"ED",X"B2",X"08",X"90",X"A7",X"CB",X"67",X"C8",
		X"96",X"09",X"9A",X"F7",X"AF",X"31",X"D8",X"27",X"89",X"0B",X"B0",X"45",X"96",X"09",X"9A",X"48",
		X"18",X"D3",X"C5",X"ED",X"B2",X"19",X"88",X"07",X"48",X"B2",X"48",X"90",X"A7",X"6F",X"46",X"01",
		X"60",X"B2",X"A8",X"38",X"87",X"EF",X"EE",X"09",X"60",X"CB",X"D0",X"C8",X"63",X"F1",X"60",X"F1",
		X"46",X"60",X"C8",X"B6",X"29",X"32",X"D7",X"87",X"31",X"F0",X"8F",X"21",X"4F",X"01",X"45",X"B6",
		X"A1",X"32",X"E0",X"38",X"F3",X"C5",X"45",X"CD",X"CD",X"80",X"65",X"BF",X"91",X"21",X"5E",X"09",
		X"CD",X"F4",X"A1",X"CD",X"54",X"29",X"21",X"1C",X"2A",X"CD",X"54",X"29",X"CD",X"F4",X"A1",X"21",
		X"15",X"0A",X"65",X"FC",X"01",X"CD",X"DC",X"81",X"89",X"51",X"A2",X"CD",X"DC",X"81",X"65",X"FC",
		X"A1",X"B6",X"D7",X"CD",X"59",X"28",X"B6",X"08",X"CD",X"46",X"3B",X"4B",X"28",X"00",X"2A",X"02",
		X"30",X"CC",X"61",X"DA",X"E5",X"CB",X"F4",X"CD",X"E4",X"80",X"E2",X"79",X"A3",X"8C",X"B0",X"EE",
		X"EF",X"CA",X"7D",X"EF",X"20",X"80",X"EB",X"EF",X"6C",X"CD",X"7A",X"49",X"2A",X"AB",X"B8",X"D8",
		X"F2",X"EF",X"E7",X"DA",X"E1",X"ED",X"E5",X"CC",X"80",X"CA",X"79",X"8B",X"25",X"98",X"E1",X"EB",
		X"E9",X"DA",X"69",X"80",X"20",X"EE",X"69",X"EB",X"69",X"EB",X"7D",X"ED",X"49",X"8A",X"3C",X"B8",
		X"E4",X"CD",X"F3",X"E9",X"E7",X"EE",X"E5",X"CC",X"80",X"CA",X"79",X"8B",X"B6",X"98",X"F3",X"E8",
		X"E9",X"EE",X"EA",X"E9",X"20",X"80",X"6D",X"CF",X"C9",X"8A",X"BE",X"98",X"6B",X"EF",X"7A",X"CD",
		X"64",X"C9",X"66",X"CC",X"80",X"DC",X"E5",X"CB",X"60",X"EE",X"67",X"EC",X"67",X"CF",X"71",X"80",
		X"E9",X"EE",X"6B",X"32",X"3A",X"80",X"3E",X"91",X"B1",X"B0",X"32",X"B2",X"B1",X"B2",X"11",X"1A",
		X"E8",X"18",X"A7",X"CE",X"E0",X"68",X"8E",X"88",X"98",X"76",X"98",X"76",X"B2",X"48",X"B8",X"07",
		X"46",X"C8",X"C8",X"1A",X"48",X"18",X"A7",X"EE",X"68",X"88",X"D0",X"89",X"A8",X"28",X"34",X"E3",
		X"2B",X"8B",X"81",X"90",X"28",X"A6",X"B0",X"6D",X"B0",X"88",X"88",X"A0",X"88",X"A0",X"88",X"A0",
		X"28",X"80",X"28",X"80",X"28",X"80",X"B2",X"48",X"18",X"0F",X"46",X"98",X"20",X"70",X"21",X"BC",
		X"28",X"94",X"81",X"A9",X"28",X"12",X"A0",X"18",X"A7",X"CE",X"27",X"30",X"12",X"81",X"91",X"28",
		X"2E",X"80",X"CD",X"98",X"28",X"80",X"28",X"80",X"28",X"80",X"28",X"80",X"28",X"80",X"28",X"80",
		X"88",X"12",X"E8",X"18",X"A7",X"CE",X"80",X"80",X"58",X"81",X"36",X"28",X"94",X"81",X"22",X"28",
		X"B2",X"88",X"18",X"0F",X"46",X"AF",X"6F",X"1A",X"28",X"18",X"A7",X"07",X"AF",X"07",X"AF",X"EE",
		X"27",X"90",X"88",X"0B",X"89",X"01",X"28",X"29",X"2B",X"0B",X"6D",X"45",X"46",X"AC",X"D9",X"0F",
		X"21",X"2D",X"2B",X"FF",X"3E",X"00",X"B9",X"FE",X"23",X"7E",X"E1",X"26",X"28",X"B9",X"45",X"F6",
		X"89",X"00",X"28",X"0E",X"DF",X"41",X"8B",X"F6",X"94",X"41",X"68",X"77",X"61",X"2D",X"A3",X"C9",
		X"2B",X"71",X"2B",X"59",X"2B",X"7C",X"2B",X"5D",X"2B",X"65",X"2B",X"52",X"2B",X"7F",X"2B",X"5F",
		X"A3",X"C4",X"A3",X"5E",X"A3",X"DF",X"A3",X"53",X"A3",X"CB",X"A3",X"45",X"A3",X"F7",X"A0",X"08",
		X"28",X"01",X"D7",X"00",X"28",X"01",X"D7",X"00",X"29",X"FF",X"29",X"FF",X"2A",X"FF",X"2B",X"FF",
		X"A4",X"F7",X"A5",X"F7",X"A6",X"F7",X"A0",X"09",X"A0",X"09",X"A1",X"09",X"5F",X"08",X"A1",X"08",
		X"2A",X"FF",X"29",X"01",X"29",X"01",X"2A",X"FF",X"29",X"01",X"29",X"02",X"D7",X"01",X"2A",X"FF",
		X"A2",X"0A",X"A2",X"0A",X"A3",X"F7",X"A2",X"0A",X"A2",X"0B",X"5F",X"2E",X"A0",X"CD",X"29",X"10",
		X"21",X"0B",X"88",X"CB",X"F6",X"C8",X"CD",X"7A",X"A3",X"21",X"1F",X"2A",X"B2",X"08",X"88",X"D6",
		X"A1",X"20",X"A3",X"21",X"08",X"82",X"65",X"FC",X"01",X"C9",X"89",X"16",X"28",X"39",X"E5",X"38",
		X"B8",X"06",X"21",X"1C",X"88",X"39",X"6C",X"90",X"F6",X"07",X"C8",X"23",X"F6",X"CB",X"F7",X"20",
		X"A6",X"36",X"2A",X"B6",X"A1",X"3A",X"61",X"46",X"57",X"A0",X"A2",X"35",X"61",X"36",X"A0",X"A3",
		X"35",X"87",X"3A",X"C9",X"21",X"00",X"18",X"2E",X"20",X"36",X"28",X"23",X"38",X"FB",X"87",X"32",
		X"E0",X"38",X"9A",X"49",X"B8",X"32",X"E3",X"38",X"9A",X"4C",X"B8",X"32",X"E5",X"38",X"9A",X"4F",
		X"18",X"32",X"6A",X"90",X"32",X"46",X"18",X"87",X"21",X"00",X"28",X"32",X"A8",X"88",X"22",X"09",
		X"28",X"92",X"23",X"28",X"82",X"BC",X"28",X"82",X"36",X"28",X"81",X"C0",X"2C",X"B1",X"C1",X"2C",
		X"29",X"FF",X"28",X"9E",X"28",X"6D",X"10",X"89",X"28",X"2F",X"39",X"89",X"8F",X"81",X"B7",X"88",
		X"96",X"88",X"65",X"98",X"6D",X"64",X"30",X"0F",X"92",X"77",X"AF",X"16",X"A1",X"92",X"E0",X"18",
		X"D3",X"2F",X"32",X"A0",X"88",X"9A",X"A1",X"28",X"21",X"88",X"28",X"8A",X"AE",X"28",X"22",X"98",
		X"28",X"81",X"F8",X"8F",X"82",X"AC",X"28",X"6D",X"E0",X"85",X"B2",X"C8",X"B8",X"07",X"8E",X"88",
		X"CB",X"D7",X"20",X"8A",X"2E",X"89",X"F0",X"9A",X"B8",X"28",X"B6",X"88",X"32",X"9F",X"88",X"89",
		X"72",X"96",X"82",X"86",X"28",X"81",X"A0",X"08",X"99",X"50",X"5F",X"8F",X"B9",X"CD",X"49",X"02",
		X"A0",X"28",X"CD",X"98",X"2D",X"9A",X"A2",X"28",X"B6",X"88",X"32",X"B9",X"88",X"65",X"00",X"8C",
		X"6D",X"81",X"A5",X"6D",X"6B",X"82",X"6D",X"41",X"A6",X"16",X"A8",X"6D",X"F9",X"A0",X"A0",X"50",
		X"B6",X"88",X"32",X"CF",X"18",X"9A",X"6A",X"18",X"32",X"CE",X"18",X"65",X"A5",X"8F",X"B8",X"78",
		X"6D",X"45",X"00",X"6D",X"9F",X"91",X"6D",X"98",X"03",X"12",X"FB",X"8C",X"76",X"80",X"48",X"81",
		X"58",X"8C",X"CD",X"54",X"A1",X"ED",X"39",X"8B",X"28",X"11",X"B6",X"80",X"96",X"E0",X"41",X"65",
		X"DC",X"A1",X"B6",X"C8",X"6D",X"59",X"00",X"6D",X"DC",X"A1",X"B6",X"48",X"6D",X"59",X"00",X"69",
		X"2A",X"AA",X"18",X"80",X"20",X"80",X"20",X"80",X"00",X"8A",X"AD",X"18",X"20",X"80",X"20",X"DC",
		X"60",X"C9",X"66",X"EB",X"F3",X"80",X"E6",X"EF",X"F2",X"80",X"F0",X"EC",X"E1",X"F9",X"61",X"EE",
		X"6F",X"B2",X"20",X"00",X"2A",X"98",X"18",X"80",X"20",X"80",X"20",X"80",X"7C",X"DA",X"F9",X"80",
		X"67",X"46",X"E3",X"4D",X"80",X"45",X"67",X"5A",X"E5",X"88",X"15",X"88",X"80",X"88",X"80",X"A8",
		X"87",X"0E",X"23",X"CB",X"6D",X"A0",X"29",X"A7",X"AB",X"FF",X"F0",X"11",X"F3",X"20",X"52",X"77",
		X"61",X"B6",X"A0",X"32",X"B6",X"20",X"65",X"ED",X"00",X"CD",X"9F",X"99",X"65",X"18",X"03",X"CD",
		X"96",X"05",X"21",X"7A",X"2D",X"45",X"39",X"03",X"28",X"B9",X"F6",X"D6",X"7B",X"20",X"42",X"41",
		X"65",X"FC",X"01",X"21",X"B8",X"0D",X"65",X"FC",X"01",X"21",X"38",X"0D",X"65",X"FC",X"01",X"26",
		X"3A",X"A6",X"2F",X"22",X"28",X"88",X"B6",X"09",X"32",X"02",X"88",X"CD",X"D6",X"2E",X"21",X"A2",
		X"A5",X"CD",X"DC",X"81",X"0E",X"1E",X"06",X"0F",X"96",X"01",X"9A",X"0A",X"28",X"CD",X"09",X"87",
		X"21",X"AE",X"2D",X"CD",X"54",X"29",X"CD",X"29",X"BD",X"C9",X"2D",X"06",X"19",X"53",X"79",X"55",
		X"E1",X"5B",X"60",X"88",X"F4",X"40",X"E5",X"88",X"F3",X"46",X"67",X"97",X"E2",X"4D",X"E5",X"7B",
		X"AC",X"0B",X"19",X"50",X"6D",X"4E",X"6F",X"CF",X"AC",X"0F",X"98",X"53",X"EE",X"4F",X"B7",X"42",
		X"E5",X"6D",X"24",X"1B",X"B9",X"41",X"E3",X"4D",X"80",X"4A",X"64",X"47",X"E3",X"63",X"24",X"1F",
		X"98",X"44",X"E9",X"41",X"ED",X"4F",X"EE",X"44",X"20",X"42",X"EC",X"4F",X"6B",X"CB",X"B6",X"09",
		X"9A",X"0A",X"28",X"B6",X"D8",X"21",X"21",X"13",X"8A",X"08",X"28",X"CD",X"A0",X"87",X"89",X"03",
		X"BB",X"22",X"28",X"88",X"CD",X"00",X"A7",X"21",X"AD",X"1B",X"22",X"00",X"88",X"CD",X"28",X"2F",
		X"89",X"07",X"33",X"22",X"A0",X"20",X"65",X"08",X"07",X"B6",X"3C",X"21",X"21",X"15",X"8A",X"08",
		X"88",X"CD",X"AC",X"06",X"B6",X"5C",X"CD",X"0C",X"2E",X"21",X"39",X"1B",X"22",X"00",X"88",X"B6",
		X"82",X"6D",X"14",X"A1",X"B4",X"6D",X"31",X"A1",X"6D",X"B4",X"01",X"69",X"8E",X"8C",X"6D",X"B4",
		X"A1",X"1C",X"38",X"72",X"C9",X"1E",X"28",X"9A",X"2A",X"28",X"21",X"D0",X"2E",X"96",X"00",X"86",
		X"20",X"ED",X"B6",X"8F",X"18",X"EE",X"A2",X"E7",X"AE",X"8D",X"65",X"E3",X"A0",X"28",X"F6",X"83",
		X"07",X"08",X"B1",X"C7",X"CB",X"5F",X"20",X"AD",X"CB",X"DF",X"20",X"9D",X"F2",X"65",X"B4",X"A1",
		X"9C",X"B0",X"59",X"30",X"49",X"CE",X"27",X"E7",X"B6",X"80",X"6D",X"B4",X"01",X"B0",X"5B",X"30",
		X"DD",X"EE",X"AF",X"ED",X"5D",X"89",X"64",X"8E",X"3E",X"88",X"FF",X"11",X"F6",X"F1",X"41",X"65",
		X"14",X"A1",X"B8",X"6A",X"8B",X"20",X"E8",X"6D",X"FB",X"44",X"48",X"61",X"49",X"B0",X"9A",X"69",
		X"2E",X"88",X"2C",X"C9",X"29",X"28",X"2B",X"88",X"2A",X"C9",X"AA",X"C8",X"2C",X"88",X"29",X"C9",
		X"A3",X"C9",X"A3",X"C9",X"E1",X"8A",X"E1",X"8C",X"A0",X"89",X"E1",X"C9",X"A1",X"C9",X"A1",X"C9",
		X"29",X"C9",X"29",X"C9",X"29",X"C9",X"2A",X"C9",X"69",X"89",X"28",X"89",X"69",X"C9",X"29",X"C9",
		X"A3",X"C9",X"A3",X"C9",X"E1",X"8A",X"E1",X"89",X"A0",X"89",X"E1",X"8A",X"E1",X"C9",X"A6",X"CB",
		X"69",X"CC",X"2A",X"88",X"29",X"CA",X"29",X"09",X"6E",X"CF",X"0C",X"8A",X"6A",X"CD",X"29",X"88",
		X"B6",X"88",X"92",X"CB",X"B8",X"6D",X"CD",X"A0",X"6D",X"17",X"91",X"6D",X"B0",X"A3",X"6D",X"E4",
		X"27",X"89",X"F6",X"8D",X"F6",X"7E",X"79",X"88",X"2E",X"1E",X"D7",X"65",X"59",X"A0",X"C9",X"E9",
		X"69",X"16",X"A5",X"92",X"B2",X"28",X"92",X"9B",X"28",X"81",X"A0",X"88",X"82",X"84",X"28",X"12",
		X"68",X"18",X"A7",X"EE",X"B8",X"07",X"AF",X"07",X"4E",X"8A",X"32",X"9C",X"88",X"9A",X"3D",X"28",
		X"A7",X"32",X"B6",X"20",X"82",X"8E",X"28",X"22",X"D8",X"24",X"89",X"52",X"96",X"22",X"86",X"20",
		X"39",X"00",X"64",X"21",X"56",X"8C",X"34",X"CB",X"6E",X"A0",X"2B",X"39",X"28",X"66",X"C5",X"7B",
		X"DA",X"24",X"A7",X"32",X"DD",X"24",X"65",X"85",X"21",X"CD",X"E8",X"0E",X"61",X"B2",X"20",X"20",
		X"07",X"C8",X"87",X"32",X"3E",X"88",X"CD",X"E5",X"A0",X"CD",X"38",X"2B",X"CD",X"2C",X"A2",X"21",
		X"23",X"20",X"63",X"D6",X"ED",X"CD",X"D4",X"0F",X"E9",X"CB",X"B6",X"B6",X"5F",X"32",X"B7",X"20",
		X"CD",X"7D",X"A8",X"87",X"32",X"17",X"88",X"32",X"6B",X"90",X"21",X"00",X"88",X"39",X"A2",X"00",
		X"AF",X"B9",X"4E",X"B2",X"02",X"20",X"B0",X"CA",X"05",X"0F",X"A7",X"A7",X"89",X"08",X"28",X"A3",
		X"77",X"4B",X"A5",X"07",X"CD",X"B7",X"31",X"DD",X"21",X"80",X"8D",X"DD",X"36",X"00",X"10",X"DD",
		X"9E",X"09",X"70",X"DD",X"9E",X"0B",X"23",X"DD",X"9E",X"0C",X"A2",X"DD",X"9E",X"0D",X"A5",X"DD",
		X"36",X"09",X"28",X"DD",X"36",X"0B",X"28",X"CD",X"CE",X"33",X"CD",X"AB",X"B1",X"CD",X"75",X"08",
		X"65",X"11",X"20",X"B2",X"A8",X"38",X"87",X"46",X"C0",X"A0",X"DA",X"CB",X"DF",X"20",X"25",X"21",
		X"A8",X"88",X"35",X"B6",X"28",X"32",X"3E",X"88",X"CD",X"D1",X"2F",X"C9",X"B2",X"08",X"88",X"D6",
		X"A1",X"A0",X"7A",X"21",X"20",X"20",X"9D",X"35",X"96",X"28",X"9A",X"1E",X"28",X"CD",X"F9",X"0F",
		X"C9",X"B2",X"28",X"90",X"A7",X"46",X"AF",X"21",X"A9",X"88",X"CD",X"FB",X"2F",X"21",X"AA",X"88",
		X"92",X"08",X"B8",X"A7",X"EE",X"07",X"4F",X"B2",X"A0",X"38",X"87",X"AF",X"07",X"AF",X"07",X"46",
		X"AF",X"90",X"20",X"03",X"21",X"09",X"88",X"CD",X"D3",X"07",X"C9",X"45",X"EE",X"0F",X"21",X"2D",
		X"A3",X"77",X"9E",X"88",X"B9",X"76",X"83",X"F6",X"E1",X"86",X"A0",X"31",X"AE",X"88",X"F6",X"9F",
		X"20",X"8C",X"AC",X"0B",X"B8",X"70",X"41",X"D9",X"C9",X"75",X"F6",X"AB",X"39",X"82",X"A8",X"E3",
		X"2F",X"A5",X"5A",X"B7",X"90",X"A8",X"74",X"A8",X"37",X"C8",X"E6",X"A8",X"74",X"A8",X"D0",X"A8",
		X"26",X"AC",X"A6",X"9B",X"22",X"88",X"88",X"65",X"28",X"A1",X"CD",X"B9",X"A1",X"1E",X"EE",X"65",
		X"14",X"A1",X"7D",X"94",X"23",X"69",X"86",X"AC",X"A6",X"9B",X"82",X"88",X"28",X"16",X"66",X"6D",
		X"B4",X"A1",X"CD",X"B9",X"A1",X"65",X"28",X"A1",X"DD",X"9C",X"AB",X"61",X"DD",X"63",X"A9",X"CE",
		X"6C",X"C7",X"20",X"6D",X"AA",X"C8",X"69",X"7D",X"96",X"AA",X"80",X"7D",X"96",X"A9",X"27",X"69",
		X"DD",X"9E",X"AB",X"88",X"C9",X"0A",X"24",X"28",X"23",X"8A",X"24",X"28",X"C9",X"89",X"28",X"88",
		X"82",X"AE",X"28",X"82",X"B0",X"28",X"B6",X"89",X"92",X"9A",X"28",X"92",X"B3",X"28",X"B2",X"C8",
		X"18",X"0F",X"46",X"B8",X"AF",X"07",X"AF",X"E6",X"2A",X"9A",X"3C",X"28",X"32",X"9D",X"88",X"89",
		X"B6",X"28",X"6B",X"56",X"80",X"A8",X"B2",X"9C",X"28",X"CE",X"57",X"68",X"B8",X"80",X"B2",X"9C",
		X"88",X"EE",X"F7",X"C7",X"B2",X"9D",X"88",X"EE",X"F7",X"47",X"08",X"60",X"CB",X"C6",X"20",X"8F",
		X"F0",X"8F",X"80",X"AA",X"94",X"30",X"DD",X"51",X"07",X"80",X"A3",X"94",X"B8",X"66",X"6D",X"F0",
		X"A0",X"65",X"5E",X"A8",X"B8",X"69",X"21",X"9E",X"88",X"63",X"F6",X"88",X"2F",X"5E",X"46",X"F7",
		X"A0",X"EB",X"B8",X"AC",X"6B",X"E6",X"4C",X"4C",X"26",X"12",X"B6",X"28",X"46",X"F6",X"A0",X"B5",
		X"CD",X"45",X"A0",X"65",X"17",X"91",X"CD",X"98",X"A3",X"65",X"76",X"A4",X"CD",X"AC",X"A5",X"65",
		X"63",X"85",X"65",X"DE",X"27",X"CD",X"75",X"86",X"65",X"DF",X"26",X"B6",X"21",X"32",X"A2",X"20",
		X"C5",X"EB",X"10",X"8D",X"CD",X"A9",X"A7",X"C5",X"EB",X"B2",X"8D",X"CD",X"81",X"2F",X"C5",X"EB",
		X"9C",X"25",X"65",X"A1",X"07",X"CD",X"C6",X"05",X"65",X"78",X"25",X"B8",X"D3",X"CD",X"2F",X"80",
		X"D6",X"11",X"20",X"03",X"B6",X"01",X"77",X"2E",X"2E",X"D6",X"2B",X"B0",X"AE",X"2E",X"A8",X"D6",
		X"20",X"B0",X"20",X"2E",X"22",X"D6",X"24",X"B0",X"A2",X"2E",X"24",X"F0",X"9A",X"68",X"2D",X"32",
		X"DD",X"8D",X"32",X"98",X"8D",X"21",X"2D",X"8D",X"39",X"20",X"28",X"36",X"29",X"B9",X"36",X"02",
		X"11",X"36",X"A3",X"B9",X"9E",X"0C",X"89",X"2D",X"2D",X"36",X"A5",X"21",X"8D",X"25",X"9E",X"0E",
		X"CD",X"E5",X"A0",X"CD",X"17",X"31",X"CD",X"10",X"A3",X"B2",X"B9",X"88",X"07",X"A0",X"2E",X"CD",
		X"D6",X"84",X"65",X"04",X"05",X"CD",X"4F",X"99",X"65",X"2B",X"92",X"CD",X"0B",X"9A",X"65",X"6A",
		X"31",X"CD",X"01",X"2D",X"B6",X"20",X"32",X"00",X"08",X"87",X"32",X"92",X"8D",X"32",X"1B",X"8D",
		X"65",X"4C",X"25",X"DD",X"89",X"28",X"2D",X"CD",X"6E",X"9B",X"65",X"A3",X"11",X"CD",X"50",X"96",
		X"CD",X"A9",X"6B",X"2E",X"D7",X"CD",X"89",X"18",X"2E",X"02",X"CD",X"89",X"B8",X"B2",X"68",X"90",
		X"87",X"CB",X"C7",X"4A",X"03",X"02",X"96",X"48",X"65",X"79",X"00",X"B2",X"C0",X"24",X"AF",X"20",
		X"D2",X"B6",X"2E",X"32",X"93",X"8C",X"87",X"21",X"FB",X"8C",X"77",X"23",X"77",X"23",X"77",X"21",
		X"7E",X"25",X"9E",X"00",X"8B",X"36",X"A8",X"B2",X"C0",X"24",X"AF",X"20",X"A7",X"53",X"0E",X"00",
		X"CD",X"89",X"B8",X"D3",X"CD",X"75",X"A8",X"CD",X"AE",X"33",X"CD",X"14",X"33",X"CD",X"BA",X"33",
		X"6D",X"80",X"93",X"6D",X"D3",X"B5",X"6D",X"36",X"E1",X"6D",X"31",X"E9",X"6D",X"AC",X"63",X"6D",
		X"E8",X"EB",X"CD",X"46",X"EB",X"65",X"7D",X"EC",X"B2",X"3E",X"8D",X"63",X"F7",X"E2",X"5A",X"AC",
		X"B2",X"38",X"2D",X"8F",X"80",X"49",X"6D",X"7D",X"23",X"10",X"1C",X"A6",X"A4",X"6D",X"29",X"B8",
		X"53",X"75",X"21",X"08",X"8D",X"1A",X"FC",X"2C",X"DD",X"A6",X"3A",X"86",X"28",X"7E",X"B4",X"18",
		X"A4",X"FE",X"14",X"A6",X"A1",X"7D",X"D7",X"9A",X"B2",X"FD",X"2C",X"7D",X"0E",X"9B",X"08",X"7D",
		X"77",X"9B",X"D3",X"65",X"B1",X"AC",X"CD",X"DD",X"AC",X"65",X"AC",X"A5",X"21",X"80",X"AB",X"65",
		X"DC",X"A1",X"81",X"B3",X"23",X"6D",X"DC",X"A1",X"81",X"DE",X"23",X"6D",X"DC",X"A1",X"81",X"D1",
		X"AB",X"65",X"54",X"A1",X"21",X"2C",X"AB",X"65",X"54",X"A1",X"21",X"07",X"AB",X"65",X"54",X"A1",
		X"81",X"4A",X"23",X"6D",X"DC",X"A1",X"B6",X"80",X"6D",X"59",X"00",X"12",X"BB",X"2D",X"86",X"88",
		X"E7",X"65",X"68",X"A3",X"26",X"8B",X"A6",X"AC",X"22",X"88",X"88",X"1E",X"38",X"9A",X"2A",X"28",
		X"6D",X"E7",X"04",X"12",X"BA",X"2D",X"86",X"88",X"E7",X"6D",X"E0",X"A3",X"86",X"8B",X"A6",X"9B",
		X"22",X"88",X"88",X"65",X"E7",X"A4",X"B6",X"80",X"CD",X"59",X"A0",X"0E",X"2A",X"8E",X"38",X"91",
		X"A0",X"88",X"7D",X"56",X"B3",X"8F",X"80",X"93",X"8E",X"89",X"6D",X"27",X"30",X"06",X"A2",X"86",
		X"AE",X"91",X"29",X"88",X"DD",X"5E",X"3A",X"7E",X"32",X"98",X"20",X"8E",X"AC",X"91",X"32",X"88",
		X"76",X"A0",X"90",X"9F",X"86",X"AA",X"99",X"C4",X"A0",X"5E",X"36",X"90",X"26",X"86",X"20",X"B1",
		X"C8",X"88",X"D6",X"9C",X"30",X"8D",X"26",X"8E",X"39",X"54",X"29",X"F5",X"B6",X"B8",X"22",X"88",
		X"28",X"2E",X"30",X"CD",X"05",X"81",X"18",X"F3",X"79",X"CD",X"0F",X"80",X"96",X"28",X"65",X"79",
		X"A0",X"CD",X"8F",X"28",X"46",X"01",X"CC",X"29",X"BD",X"CD",X"8F",X"28",X"34",X"4B",X"A5",X"09",
		X"A2",X"0B",X"30",X"4F",X"E1",X"45",X"E5",X"88",X"F4",X"41",X"65",X"4D",X"80",X"88",X"80",X"88",
		X"ED",X"49",X"EE",X"3A",X"20",X"20",X"20",X"53",X"6D",X"43",X"92",X"02",X"2E",X"11",X"6E",X"52",
		X"67",X"45",X"80",X"98",X"90",X"88",X"F4",X"47",X"80",X"99",X"11",X"88",X"12",X"9D",X"90",X"98",
		X"30",X"20",X"78",X"54",X"7B",X"BA",X"2A",X"08",X"39",X"46",X"7A",X"4F",X"ED",X"20",X"32",X"30",
		X"80",X"5C",X"67",X"88",X"92",X"91",X"80",X"92",X"92",X"98",X"90",X"98",X"80",X"58",X"F4",X"5B",
		X"92",X"02",X"AA",X"11",X"6E",X"52",X"EF",X"4D",X"20",X"33",X"30",X"20",X"7C",X"4F",X"20",X"33",
		X"11",X"88",X"12",X"99",X"90",X"98",X"90",X"88",X"F0",X"5C",X"F3",X"B2",X"A2",X"04",X"B1",X"4E",
		X"7A",X"4F",X"ED",X"20",X"34",X"30",X"20",X"54",X"EF",X"20",X"34",X"39",X"20",X"3A",X"B2",X"35",
		X"90",X"98",X"80",X"58",X"F4",X"5B",X"1A",X"0A",X"26",X"19",X"E6",X"5A",X"67",X"45",X"80",X"9D",
		X"30",X"20",X"7C",X"4F",X"20",X"35",X"B1",X"20",X"B2",X"3A",X"B2",X"31",X"30",X"20",X"78",X"54",
		X"F3",X"B2",X"A2",X"18",X"B1",X"9E",X"90",X"88",X"E1",X"46",X"E4",X"88",X"67",X"5E",X"E5",X"5A",
		X"20",X"20",X"20",X"20",X"EE",X"4F",X"20",X"42",X"EF",X"4E",X"7D",X"53",X"92",X"CD",X"C4",X"0B",
		X"65",X"F1",X"23",X"D8",X"65",X"16",X"24",X"D8",X"65",X"8E",X"24",X"C9",X"89",X"37",X"2D",X"F6",
		X"D6",X"02",X"B0",X"04",X"20",X"02",X"36",X"01",X"C9",X"21",X"BF",X"8D",X"39",X"20",X"28",X"2E",
		X"A4",X"56",X"76",X"8A",X"B0",X"8C",X"80",X"8A",X"96",X"89",X"B9",X"B0",X"DC",X"81",X"37",X"2D",
		X"2E",X"8C",X"F6",X"7E",X"2B",X"18",X"2A",X"9F",X"C9",X"11",X"38",X"56",X"07",X"61",X"21",X"37",
		X"2D",X"56",X"07",X"68",X"97",X"69",X"81",X"4D",X"2C",X"B1",X"A6",X"88",X"8E",X"8C",X"F6",X"8F",
		X"20",X"8D",X"B9",X"90",X"D1",X"AF",X"C9",X"9F",X"C9",X"86",X"20",X"E5",X"B6",X"80",X"18",X"1C",
		X"CF",X"26",X"A0",X"4D",X"CB",X"88",X"28",X"16",X"A0",X"6D",X"90",X"A7",X"B6",X"89",X"6D",X"59",
		X"A0",X"E1",X"38",X"47",X"C9",X"75",X"21",X"08",X"8D",X"75",X"F6",X"88",X"DD",X"9E",X"2C",X"8A",
		X"76",X"08",X"90",X"8C",X"7D",X"96",X"A4",X"8B",X"7D",X"96",X"A6",X"AF",X"7D",X"96",X"20",X"77",
		X"CD",X"D5",X"A8",X"86",X"08",X"90",X"D6",X"65",X"EA",X"B1",X"DD",X"9C",X"2F",X"75",X"F6",X"8F",
		X"7D",X"1E",X"A6",X"10",X"4B",X"7D",X"96",X"8F",X"A0",X"7D",X"F6",X"88",X"07",X"68",X"76",X"68",
		X"CC",X"00",X"AC",X"75",X"F6",X"88",X"D6",X"A0",X"CC",X"31",X"AC",X"65",X"5F",X"B5",X"B8",X"58",
		X"7D",X"56",X"A4",X"5E",X"A3",X"E8",X"6D",X"F4",X"05",X"CE",X"A1",X"68",X"7D",X"96",X"A2",X"40",
		X"CD",X"23",X"B1",X"1E",X"68",X"65",X"59",X"A0",X"C9",X"75",X"F6",X"8C",X"D6",X"8A",X"48",X"65",
		X"54",X"A5",X"46",X"89",X"68",X"7D",X"96",X"8A",X"CA",X"6D",X"0B",X"B1",X"B6",X"C8",X"6D",X"59",
		X"A0",X"61",X"CD",X"40",X"AB",X"72",X"47",X"A9",X"2E",X"8D",X"CD",X"29",X"B8",X"1E",X"2E",X"9A",
		X"3F",X"2D",X"7D",X"81",X"A8",X"2D",X"6D",X"13",X"17",X"16",X"A6",X"7D",X"36",X"BF",X"A0",X"52",
		X"53",X"75",X"21",X"08",X"8D",X"1A",X"FC",X"2C",X"DD",X"A6",X"3A",X"86",X"28",X"7E",X"B4",X"18",
		X"A4",X"5E",X"14",X"2E",X"A1",X"DD",X"DF",X"1A",X"92",X"55",X"2C",X"DD",X"2E",X"1B",X"28",X"DD",
		X"77",X"13",X"D3",X"B6",X"28",X"32",X"9E",X"8D",X"CD",X"9E",X"A0",X"F6",X"B5",X"77",X"46",X"7F",
		X"62",X"7F",X"26",X"B2",X"31",X"20",X"AF",X"C8",X"96",X"28",X"65",X"79",X"00",X"CD",X"11",X"04",
		X"CD",X"38",X"AE",X"21",X"3E",X"88",X"CB",X"F6",X"A0",X"07",X"34",X"CB",X"6E",X"CC",X"4C",X"0E",
		X"61",X"34",X"9C",X"C9",X"65",X"36",X"00",X"D6",X"A5",X"58",X"95",X"0F",X"8E",X"8B",X"C7",X"22",
		X"28",X"88",X"45",X"CD",X"28",X"29",X"CD",X"00",X"A1",X"41",X"26",X"00",X"22",X"00",X"88",X"CD",
		X"A0",X"81",X"65",X"08",X"01",X"C9",X"75",X"21",X"A8",X"25",X"89",X"35",X"25",X"EE",X"8B",X"6E",
		X"23",X"45",X"CD",X"0A",X"30",X"B0",X"23",X"CD",X"87",X"0D",X"B0",X"1E",X"41",X"F1",X"4E",X"02",
		X"2F",X"0F",X"2F",X"DD",X"DF",X"08",X"D0",X"0F",X"2F",X"0F",X"75",X"77",X"A1",X"DD",X"9E",X"0A",
		X"A8",X"DD",X"36",X"1E",X"28",X"DD",X"36",X"1F",X"29",X"C9",X"41",X"B8",X"58",X"0D",X"AE",X"0D",
		X"24",X"05",X"B0",X"03",X"26",X"07",X"26",X"03",X"B0",X"07",X"B0",X"03",X"24",X"07",X"24",X"4D",
		X"78",X"F9",X"A2",X"B0",X"8D",X"CD",X"99",X"2D",X"A0",X"13",X"A2",X"B2",X"8D",X"CD",X"99",X"2D",
		X"80",X"03",X"82",X"BC",X"2D",X"CD",X"39",X"85",X"80",X"0B",X"69",X"87",X"61",X"49",X"9F",X"C9",
		X"21",X"2C",X"AE",X"DD",X"21",X"00",X"8D",X"DD",X"F6",X"1F",X"07",X"4C",X"28",X"0E",X"DD",X"21",
		X"80",X"25",X"75",X"F6",X"37",X"07",X"6C",X"08",X"26",X"DD",X"89",X"48",X"2D",X"DD",X"D6",X"17",
		X"07",X"4C",X"28",X"0E",X"DD",X"21",X"60",X"8D",X"DD",X"F6",X"BF",X"07",X"4C",X"00",X"AE",X"C9",
		X"EE",X"83",X"CE",X"83",X"DE",X"83",X"45",X"FD",X"6D",X"E7",X"01",X"16",X"80",X"1E",X"A0",X"8E",
		X"59",X"58",X"0A",X"C7",X"B8",X"51",X"59",X"59",X"4E",X"8A",X"0F",X"A7",X"0F",X"75",X"77",X"88",
		X"F0",X"AF",X"0F",X"AF",X"7D",X"D7",X"A1",X"6D",X"6E",X"93",X"41",X"69",X"A1",X"8A",X"A2",X"B9",
		X"BE",X"76",X"B9",X"8A",X"2A",X"89",X"BE",X"76",X"21",X"40",X"8D",X"86",X"2A",X"E5",X"AE",X"AD",
		X"4D",X"16",X"A2",X"B8",X"0F",X"AF",X"0F",X"AF",X"4E",X"8A",X"DF",X"16",X"25",X"B9",X"0F",X"EE",
		X"29",X"57",X"CD",X"FD",X"AE",X"E1",X"AD",X"88",X"47",X"E1",X"38",X"41",X"C9",X"9E",X"28",X"86",
		X"20",X"ED",X"5D",X"E2",X"EB",X"CD",X"6D",X"E7",X"01",X"56",X"41",X"5E",X"80",X"6B",X"9E",X"F9",
		X"49",X"94",X"3C",X"90",X"C4",X"8B",X"C9",X"1E",X"28",X"9A",X"2A",X"28",X"21",X"40",X"8D",X"86",
		X"A2",X"ED",X"AE",X"AD",X"4D",X"16",X"25",X"B9",X"0F",X"EE",X"A1",X"77",X"F0",X"B6",X"A2",X"15",
		X"A0",X"8D",X"CD",X"23",X"AE",X"10",X"2D",X"96",X"3A",X"65",X"07",X"AE",X"49",X"05",X"20",X"44",
		X"49",X"B0",X"7E",X"6D",X"B4",X"A7",X"69",X"A6",X"A7",X"30",X"A2",X"A6",X"20",X"ED",X"5D",X"4D",
		X"7B",X"88",X"88",X"63",X"3E",X"98",X"2D",X"ED",X"CD",X"76",X"A6",X"E9",X"59",X"E1",X"3C",X"94",
		X"98",X"63",X"83",X"69",X"81",X"88",X"2D",X"B1",X"A0",X"2E",X"8E",X"88",X"F6",X"DD",X"BA",X"D7",
		X"51",X"92",X"23",X"93",X"38",X"56",X"C9",X"65",X"17",X"91",X"2E",X"8E",X"CD",X"29",X"B8",X"89",
		X"64",X"AF",X"6D",X"A6",X"27",X"81",X"F1",X"AF",X"B2",X"9E",X"28",X"6B",X"CF",X"00",X"A3",X"81",
		X"FD",X"AF",X"CD",X"54",X"A1",X"89",X"E1",X"AF",X"CD",X"54",X"A1",X"1E",X"08",X"65",X"59",X"A0",
		X"65",X"27",X"85",X"21",X"B6",X"20",X"63",X"F6",X"80",X"0F",X"9C",X"CB",X"4E",X"CC",X"EC",X"06",
		X"C9",X"34",X"34",X"21",X"28",X"84",X"3E",X"04",X"BE",X"2A",X"B9",X"EE",X"21",X"00",X"08",X"3E",
		X"5F",X"BE",X"D8",X"B9",X"D6",X"91",X"60",X"21",X"A0",X"20",X"83",X"36",X"5F",X"C9",X"56",X"23",
		X"7E",X"23",X"F6",X"32",X"2A",X"88",X"23",X"EE",X"23",X"6E",X"4D",X"5D",X"C5",X"7B",X"28",X"88",
		X"65",X"08",X"01",X"AD",X"88",X"F2",X"79",X"49",X"1C",X"38",X"4F",X"C9",X"20",X"04",X"B0",X"04",
		X"2D",X"09",X"AD",X"10",X"78",X"4C",X"69",X"59",X"6D",X"52",X"20",X"20",X"11",X"09",X"AD",X"10",
		X"F0",X"44",X"E1",X"51",X"E5",X"5A",X"80",X"88",X"9A",X"01",X"27",X"18",X"E7",X"49",X"65",X"4D",
		X"20",X"20",X"EF",X"56",X"6D",X"D2",X"21",X"E3",X"AF",X"B2",X"3E",X"88",X"CB",X"6F",X"A0",X"03",
		X"89",X"E6",X"27",X"CD",X"DC",X"81",X"89",X"F1",X"27",X"CD",X"DC",X"81",X"96",X"28",X"65",X"79",
		X"A0",X"21",X"DE",X"0F",X"CD",X"2E",X"AF",X"C9",X"2E",X"10",X"AE",X"09",X"3E",X"05",X"BE",X"0A",
		X"89",X"8F",X"2C",X"5D",X"6D",X"5D",X"ED",X"CD",X"47",X"81",X"D6",X"41",X"DF",X"23",X"04",X"59",
		X"BD",X"20",X"52",X"49",X"2C",X"59",X"3D",X"20",X"C2",X"C9",X"2E",X"10",X"AE",X"09",X"3E",X"05",
		X"16",X"02",X"89",X"8F",X"2C",X"5D",X"6D",X"5D",X"ED",X"F6",X"FD",X"CD",X"47",X"81",X"F9",X"77",
		X"41",X"23",X"AC",X"59",X"BD",X"20",X"50",X"49",X"2C",X"59",X"3D",X"20",X"C0",X"C9",X"A9",X"10",
		X"A0",X"02",X"A5",X"02",X"B1",X"18",X"F0",X"44",X"E1",X"51",X"E5",X"5A",X"80",X"B9",X"22",X"19",
		X"38",X"50",X"EC",X"41",X"F9",X"45",X"7A",X"20",X"12",X"0B",X"3B",X"10",X"7A",X"45",X"69",X"44",
		X"D9",X"FF",X"D7",X"B6",X"28",X"BA",X"6F",X"90",X"BA",X"42",X"18",X"BA",X"6E",X"90",X"45",X"F2",
		X"10",X"6D",X"BF",X"31",X"65",X"69",X"90",X"6D",X"1B",X"38",X"65",X"3C",X"93",X"6D",X"1B",X"38",
		X"45",X"F1",X"3C",X"45",X"B3",X"10",X"45",X"66",X"3C",X"45",X"B3",X"10",X"45",X"0D",X"39",X"45",
		X"1B",X"38",X"65",X"76",X"96",X"6D",X"1B",X"38",X"E3",X"28",X"80",X"B6",X"02",X"6D",X"F1",X"A0",
		X"41",X"55",X"CB",X"26",X"28",X"A9",X"28",X"80",X"45",X"F2",X"38",X"B0",X"2A",X"43",X"49",X"A9",
		X"80",X"88",X"65",X"52",X"90",X"B0",X"82",X"6B",X"61",X"7D",X"EB",X"6D",X"ED",X"A0",X"89",X"09",
		X"38",X"45",X"54",X"29",X"45",X"D2",X"38",X"45",X"42",X"10",X"A9",X"8F",X"38",X"F1",X"8F",X"A0",
		X"83",X"81",X"35",X"38",X"FD",X"6D",X"FC",X"A1",X"F9",X"80",X"7E",X"B6",X"82",X"6D",X"C6",X"3B",
		X"41",X"08",X"AA",X"10",X"7A",X"41",X"ED",X"53",X"20",X"20",X"20",X"54",X"6D",X"53",X"5C",X"08",
		X"92",X"38",X"C1",X"EC",X"44",X"20",X"D2",X"69",X"45",X"7B",X"88",X"EF",X"63",X"A8",X"92",X"3E",
		X"7A",X"41",X"ED",X"53",X"20",X"42",X"69",X"C4",X"A8",X"0D",X"38",X"52",X"69",X"4D",X"31",X"20",
		X"47",X"CB",X"00",X"AD",X"96",X"7A",X"C1",X"ED",X"99",X"20",X"C2",X"69",X"E4",X"A8",X"07",X"38",
		X"7A",X"41",X"ED",X"32",X"20",X"4F",X"CB",X"08",X"AF",X"16",X"7A",X"41",X"ED",X"32",X"20",X"42",
		X"C1",X"4C",X"89",X"80",X"90",X"6B",X"C1",X"A0",X"83",X"81",X"BA",X"38",X"E5",X"6D",X"FC",X"A1",
		X"49",X"41",X"A9",X"BD",X"38",X"43",X"61",X"A0",X"2B",X"A9",X"4F",X"10",X"4D",X"45",X"54",X"29",
		X"E1",X"69",X"7D",X"43",X"D1",X"89",X"80",X"A8",X"1E",X"7D",X"DF",X"36",X"E0",X"B6",X"2A",X"D7",
		X"B6",X"C0",X"8B",X"0B",X"D0",X"B1",X"80",X"D8",X"42",X"FD",X"EB",X"AF",X"61",X"CD",X"CD",X"A0",
		X"89",X"BE",X"92",X"65",X"FC",X"A1",X"89",X"A5",X"92",X"65",X"FC",X"A1",X"89",X"B7",X"92",X"65",
		X"DC",X"A1",X"92",X"68",X"18",X"CD",X"42",X"39",X"89",X"6E",X"3A",X"CD",X"DC",X"A1",X"92",X"28",
		X"B0",X"65",X"62",X"39",X"89",X"ED",X"92",X"65",X"FC",X"A1",X"1A",X"68",X"B0",X"87",X"63",X"47",
		X"88",X"2E",X"89",X"76",X"3A",X"CD",X"DC",X"A1",X"89",X"EC",X"3A",X"3A",X"68",X"18",X"87",X"CB",
		X"D7",X"80",X"83",X"89",X"D9",X"3A",X"65",X"54",X"09",X"92",X"C0",X"18",X"0F",X"07",X"07",X"07",
		X"EE",X"2B",X"6E",X"2A",X"FE",X"B8",X"89",X"2C",X"3B",X"22",X"28",X"00",X"65",X"B4",X"A1",X"21",
		X"5C",X"3A",X"65",X"54",X"09",X"89",X"A6",X"3A",X"65",X"54",X"09",X"92",X"C0",X"18",X"0F",X"63",
		X"C7",X"20",X"2E",X"21",X"1D",X"3A",X"65",X"DC",X"A1",X"21",X"13",X"3A",X"65",X"DC",X"A1",X"3A",
		X"C0",X"18",X"0F",X"63",X"DF",X"80",X"86",X"89",X"2E",X"3A",X"65",X"54",X"09",X"89",X"EE",X"3A",
		X"92",X"68",X"18",X"2F",X"0F",X"07",X"EE",X"2B",X"80",X"39",X"89",X"C5",X"3A",X"FE",X"29",X"28",
		X"02",X"89",X"FE",X"3A",X"7E",X"2A",X"08",X"2B",X"89",X"D5",X"92",X"65",X"FC",X"A1",X"89",X"2F",
		X"3B",X"CD",X"DC",X"A1",X"96",X"36",X"65",X"6E",X"3B",X"C9",X"87",X"06",X"20",X"0E",X"67",X"0F",
		X"98",X"2A",X"06",X"6B",X"FD",X"D1",X"65",X"B4",X"09",X"65",X"80",X"A1",X"F9",X"18",X"6E",X"61",
		X"EE",X"27",X"2F",X"16",X"28",X"5F",X"89",X"D6",X"39",X"19",X"96",X"22",X"9A",X"28",X"00",X"7E",
		X"65",X"B4",X"09",X"8B",X"1E",X"39",X"9A",X"28",X"20",X"D6",X"65",X"B4",X"09",X"61",X"9C",X"31",
		X"33",X"31",X"32",X"31",X"31",X"31",X"31",X"32",X"31",X"33",X"31",X"34",X"31",X"35",X"31",X"36",
		X"45",X"6A",X"45",X"6A",X"45",X"6A",X"45",X"6A",X"45",X"6A",X"45",X"6A",X"45",X"6A",X"00",X"2C",
		X"38",X"44",X"E9",X"50",X"20",X"53",X"7F",X"49",X"7C",X"43",X"E8",X"45",X"5B",X"08",X"2E",X"10",
		X"99",X"20",X"9A",X"20",X"9B",X"20",X"9C",X"20",X"9D",X"20",X"9E",X"20",X"9F",X"20",X"38",X"2C",
		X"A8",X"10",X"31",X"53",X"7F",X"A0",X"2C",X"0A",X"38",X"32",X"7B",X"57",X"00",X"04",X"AF",X"18",
		X"C4",X"6D",X"45",X"EF",X"88",X"7B",X"47",X"7D",X"46",X"6C",X"D3",X"20",X"47",X"CE",X"90",X"AF",
		X"B8",X"4F",X"6E",X"C6",X"2C",X"11",X"38",X"54",X"69",X"42",X"EC",X"45",X"20",X"54",X"F9",X"50",
		X"E5",X"2C",X"91",X"38",X"D5",X"78",X"88",X"7A",X"41",X"6F",X"40",X"5C",X"86",X"3B",X"10",X"78",
		X"6D",X"4E",X"6F",X"4F",X"6D",X"D3",X"2C",X"15",X"38",X"52",X"69",X"43",X"EB",X"20",X"7C",X"45",
		X"D3",X"7C",X"88",X"EF",X"66",X"AE",X"95",X"38",X"47",X"6E",X"E6",X"2C",X"05",X"38",X"C2",X"EF",
		X"EE",X"55",X"7B",X"20",X"35",X"30",X"30",X"30",X"30",X"20",X"78",X"54",X"7B",X"BA",X"AA",X"0D",
		X"90",X"33",X"98",X"30",X"98",X"10",X"84",X"B9",X"90",X"6B",X"47",X"E9",X"46",X"31",X"88",X"20",
		X"20",X"43",X"EF",X"49",X"EE",X"20",X"20",X"20",X"6B",X"52",X"6D",X"44",X"E9",X"D4",X"2C",X"1B",
		X"90",X"6B",X"47",X"E9",X"46",X"32",X"88",X"20",X"88",X"6B",X"47",X"E9",X"46",X"20",X"88",X"20",
		X"6B",X"52",X"6D",X"44",X"E9",X"D4",X"AF",X"17",X"B8",X"45",X"69",X"53",X"D9",X"0F",X"3F",X"18",
		X"45",X"6D",X"C4",X"E9",X"D5",X"CD",X"07",X"3F",X"10",X"E8",X"C1",X"7A",X"E4",X"AF",X"97",X"B8",
		X"60",X"69",X"7A",X"6C",X"6D",X"7B",X"5C",X"2C",X"3F",X"30",X"6C",X"61",X"6E",X"6E",X"61",X"6B",
		X"D5",X"EC",X"D4",X"D9",X"65",X"45",X"08",X"89",X"CC",X"3B",X"65",X"54",X"09",X"A7",X"9A",X"60",
		X"00",X"CD",X"57",X"3B",X"65",X"D6",X"3B",X"CD",X"35",X"3C",X"65",X"B4",X"3C",X"21",X"FA",X"3B",
		X"1A",X"60",X"20",X"AF",X"08",X"2B",X"89",X"08",X"93",X"FD",X"65",X"54",X"09",X"F9",X"88",X"D6",
		X"96",X"2A",X"65",X"6E",X"3B",X"C9",X"4F",X"C5",X"65",X"78",X"3B",X"C1",X"70",X"10",X"D0",X"C9",
		X"86",X"68",X"E5",X"96",X"81",X"65",X"F1",X"A0",X"E1",X"92",X"A0",X"18",X"63",X"C7",X"9F",X"60",
		X"18",X"D8",X"AF",X"C9",X"20",X"22",X"38",X"6D",X"78",X"7A",X"67",X"65",X"7B",X"A8",X"7C",X"6D",
		X"D3",X"5C",X"00",X"B8",X"90",X"69",X"44",X"EC",X"88",X"7A",X"47",X"ED",X"D3",X"20",X"47",X"CB",
		X"20",X"30",X"3E",X"6A",X"69",X"6C",X"A8",X"7A",X"67",X"65",X"5B",X"20",X"26",X"38",X"7A",X"67",
		X"45",X"31",X"88",X"EF",X"63",X"A8",X"06",X"3E",X"D2",X"EF",X"45",X"31",X"88",X"6A",X"C1",X"4C",
		X"20",X"38",X"38",X"7A",X"67",X"65",X"BA",X"A8",X"67",X"43",X"20",X"38",X"3E",X"7A",X"67",X"65",
		X"9A",X"20",X"C2",X"69",X"E4",X"A8",X"92",X"38",X"D2",X"EF",X"45",X"33",X"88",X"EF",X"63",X"A8",
		X"3A",X"3E",X"7A",X"67",X"65",X"BB",X"A8",X"6A",X"69",X"4C",X"20",X"3C",X"38",X"7A",X"67",X"65",
		X"9C",X"20",X"47",X"CB",X"00",X"3C",X"96",X"7A",X"47",X"ED",X"9C",X"20",X"C2",X"69",X"E4",X"89",
		X"28",X"28",X"09",X"28",X"A8",X"CD",X"73",X"3C",X"89",X"D0",X"F7",X"77",X"B6",X"21",X"03",X"3B",
		X"08",X"A8",X"1E",X"D7",X"9A",X"60",X"20",X"89",X"B5",X"3B",X"65",X"54",X"09",X"61",X"89",X"28",
		X"20",X"29",X"28",X"20",X"45",X"5B",X"3C",X"A9",X"D2",X"7F",X"FF",X"96",X"A9",X"A0",X"3B",X"A0",
		X"00",X"B6",X"7F",X"92",X"C8",X"88",X"89",X"82",X"93",X"6D",X"FC",X"A1",X"61",X"81",X"80",X"68",
		X"29",X"00",X"20",X"45",X"FB",X"14",X"A9",X"FC",X"F7",X"FF",X"96",X"A9",X"15",X"13",X"A0",X"08",
		X"1E",X"D7",X"9A",X"60",X"20",X"81",X"3F",X"3B",X"65",X"54",X"09",X"69",X"89",X"28",X"C8",X"89",
		X"D0",X"1F",X"45",X"5B",X"3C",X"A9",X"D6",X"7F",X"FF",X"96",X"A9",X"CA",X"3B",X"A0",X"A8",X"B6",
		X"7F",X"92",X"C8",X"88",X"89",X"5C",X"93",X"6D",X"FC",X"A1",X"61",X"27",X"A6",X"83",X"03",X"DF",
		X"F0",X"99",X"F2",X"A8",X"57",X"41",X"45",X"E5",X"A0",X"A9",X"28",X"00",X"AA",X"00",X"88",X"45",
		X"E6",X"3C",X"89",X"BB",X"80",X"82",X"80",X"88",X"65",X"4E",X"94",X"81",X"80",X"22",X"8A",X"28",
		X"88",X"45",X"D8",X"14",X"A9",X"00",X"3C",X"AA",X"28",X"88",X"45",X"D8",X"3C",X"A9",X"28",X"21",
		X"8A",X"28",X"20",X"6D",X"70",X"3C",X"89",X"2B",X"06",X"82",X"80",X"88",X"1E",X"3B",X"9A",X"2A",
		X"88",X"45",X"47",X"14",X"A9",X"03",X"38",X"AA",X"28",X"88",X"B6",X"17",X"BA",X"02",X"88",X"45",
		X"EF",X"3C",X"89",X"2B",X"92",X"82",X"80",X"88",X"1E",X"3E",X"9A",X"2A",X"20",X"6D",X"EF",X"3C",
		X"B6",X"3C",X"45",X"46",X"3B",X"41",X"2E",X"24",X"B6",X"10",X"BA",X"02",X"88",X"B6",X"2B",X"45",
		X"1C",X"A1",X"65",X"B9",X"09",X"98",X"78",X"69",X"86",X"BC",X"1E",X"38",X"9A",X"2A",X"20",X"B6",
		X"2B",X"45",X"B4",X"29",X"38",X"FB",X"41",X"2E",X"3E",X"B6",X"2B",X"45",X"B4",X"29",X"38",X"FB",
		X"61",X"6D",X"ED",X"A0",X"1E",X"38",X"9A",X"2A",X"20",X"81",X"53",X"3E",X"91",X"2E",X"84",X"65",
		X"5B",X"28",X"00",X"CD",X"4E",X"3D",X"19",X"2E",X"2F",X"ED",X"5B",X"28",X"00",X"CD",X"4E",X"3D",
		X"91",X"A9",X"02",X"65",X"EB",X"3D",X"1A",X"68",X"B0",X"EE",X"84",X"80",X"10",X"19",X"01",X"39",
		X"65",X"CB",X"3D",X"21",X"7F",X"3E",X"19",X"2E",X"22",X"CD",X"5C",X"3D",X"89",X"71",X"3E",X"11",
		X"86",X"39",X"65",X"5C",X"95",X"19",X"88",X"2A",X"86",X"AA",X"06",X"D7",X"1A",X"08",X"B0",X"89",
		X"32",X"3E",X"EE",X"A8",X"88",X"20",X"B3",X"28",X"2A",X"15",X"60",X"21",X"37",X"3E",X"57",X"C5",
		X"F5",X"19",X"01",X"2F",X"6D",X"5B",X"80",X"88",X"65",X"4E",X"95",X"92",X"A0",X"18",X"89",X"BA",
		X"3E",X"E6",X"68",X"20",X"2B",X"21",X"37",X"3E",X"19",X"3B",X"2F",X"ED",X"5B",X"28",X"00",X"CD",
		X"E6",X"3D",X"1A",X"48",X"B0",X"19",X"92",X"AA",X"65",X"98",X"95",X"92",X"C0",X"18",X"EE",X"2C",
		X"80",X"21",X"92",X"08",X"18",X"11",X"3A",X"39",X"65",X"10",X"3D",X"3E",X"29",X"CD",X"59",X"A0",
		X"F1",X"69",X"05",X"88",X"AF",X"18",X"AD",X"61",X"81",X"29",X"84",X"FD",X"89",X"24",X"96",X"A9",
		X"80",X"2B",X"89",X"AF",X"3E",X"ED",X"5B",X"28",X"00",X"C5",X"65",X"4E",X"3D",X"C1",X"F9",X"14",
		X"63",X"09",X"90",X"47",X"89",X"24",X"96",X"EE",X"A0",X"80",X"83",X"89",X"8F",X"3E",X"6D",X"5B",
		X"28",X"00",X"65",X"4E",X"3D",X"C9",X"D6",X"23",X"47",X"E6",X"F7",X"CD",X"B4",X"A1",X"D1",X"E6",
		X"A0",X"80",X"FB",X"61",X"86",X"2D",X"ED",X"E5",X"D3",X"28",X"20",X"65",X"E6",X"3D",X"E9",X"1C",
		X"18",X"DC",X"61",X"21",X"A2",X"3E",X"E5",X"53",X"28",X"00",X"1C",X"CD",X"4E",X"3D",X"89",X"BB",
		X"96",X"E5",X"D3",X"28",X"20",X"1C",X"65",X"4E",X"95",X"89",X"1C",X"3E",X"6D",X"5B",X"80",X"88",
		X"3C",X"45",X"4E",X"15",X"A9",X"45",X"3E",X"C5",X"7B",X"00",X"88",X"3C",X"45",X"C6",X"3D",X"A9",
		X"46",X"3E",X"6D",X"DB",X"80",X"88",X"65",X"4E",X"95",X"69",X"88",X"20",X"88",X"20",X"A8",X"7B",
		X"7C",X"41",X"7A",X"D4",X"20",X"4F",X"CE",X"4F",X"6E",X"C6",X"7D",X"50",X"B2",X"3A",X"B2",X"3A",
		X"1A",X"B2",X"3A",X"6C",X"47",X"7F",X"46",X"B2",X"1A",X"B2",X"1A",X"92",X"44",X"6D",X"C6",X"7C",
		X"B2",X"3A",X"B2",X"3A",X"92",X"52",X"E9",X"47",X"E8",X"54",X"B2",X"3A",X"B2",X"BA",X"78",X"55",
		X"D3",X"E8",X"1A",X"B2",X"1A",X"B2",X"3A",X"78",X"B9",X"78",X"BA",X"78",X"44",X"69",X"51",X"6D",
		X"7A",X"20",X"6B",X"4F",X"EE",X"54",X"7A",X"4F",X"EC",X"D3",X"31",X"50",X"20",X"20",X"20",X"20",
		X"88",X"20",X"88",X"20",X"9A",X"58",X"FB",X"B6",X"84",X"92",X"83",X"8C",X"65",X"10",X"96",X"B6",
		X"B4",X"45",X"DF",X"16",X"A0",X"28",X"F0",X"8F",X"42",X"AE",X"3E",X"BA",X"28",X"8C",X"45",X"16",
		X"97",X"8E",X"80",X"7A",X"A9",X"3E",X"65",X"09",X"97",X"8E",X"81",X"5A",X"A9",X"3E",X"65",X"94",
		X"3F",X"45",X"9B",X"17",X"A9",X"03",X"8C",X"BC",X"B6",X"20",X"96",X"4A",X"F7",X"16",X"D3",X"41",
		X"65",X"45",X"08",X"81",X"E0",X"3E",X"65",X"54",X"09",X"81",X"65",X"3E",X"65",X"54",X"09",X"69",
		X"A8",X"00",X"38",X"43",X"EF",X"49",X"EE",X"53",X"20",X"54",X"6D",X"53",X"5C",X"06",X"2A",X"10",
		X"C2",X"69",X"C4",X"20",X"88",X"20",X"C7",X"EF",X"47",X"6C",X"88",X"20",X"C2",X"69",X"E4",X"DF",
		X"5D",X"45",X"C2",X"16",X"59",X"48",X"3D",X"A8",X"57",X"41",X"3E",X"65",X"36",X"00",X"45",X"F8",
		X"96",X"48",X"13",X"F2",X"AF",X"80",X"FF",X"69",X"86",X"28",X"1A",X"08",X"B0",X"A7",X"63",X"E7",
		X"68",X"3A",X"48",X"18",X"0E",X"69",X"87",X"CB",X"CF",X"C0",X"0C",X"3A",X"48",X"18",X"87",X"CB",
		X"4F",X"68",X"9A",X"70",X"B0",X"61",X"1E",X"2D",X"9A",X"2A",X"24",X"96",X"8C",X"9A",X"81",X"8C",
		X"65",X"72",X"3F",X"CD",X"EF",X"3F",X"92",X"2A",X"04",X"90",X"9A",X"2A",X"04",X"CD",X"72",X"3F",
		X"65",X"67",X"97",X"D0",X"AF",X"62",X"41",X"3F",X"89",X"29",X"24",X"9D",X"89",X"2A",X"24",X"9D",
		X"62",X"61",X"3F",X"CD",X"72",X"3F",X"6B",X"B8",X"3F",X"CD",X"72",X"3F",X"89",X"29",X"04",X"35",
		X"E2",X"E9",X"97",X"92",X"82",X"8C",X"AF",X"60",X"9F",X"61",X"86",X"2C",X"06",X"93",X"05",X"88",
		X"D5",X"10",X"D1",X"32",X"F8",X"18",X"61",X"06",X"28",X"3A",X"28",X"04",X"F6",X"69",X"6A",X"F1",
		X"97",X"92",X"E0",X"18",X"63",X"CF",X"E0",X"0C",X"61",X"92",X"E0",X"18",X"63",X"C7",X"E0",X"0C",
		X"61",X"3E",X"AC",X"32",X"29",X"04",X"65",X"72",X"3F",X"CD",X"EF",X"3F",X"D0",X"A7",X"62",X"1B",
		X"97",X"9F",X"61",X"89",X"81",X"8C",X"9D",X"6A",X"A6",X"3F",X"61",X"D0",X"86",X"2F",X"AF",X"62",
		X"83",X"3F",X"0E",X"25",X"F6",X"29",X"62",X"83",X"3F",X"06",X"3B",X"78",X"9A",X"28",X"00",X"3A",
		X"83",X"8C",X"9A",X"29",X"20",X"92",X"80",X"8C",X"65",X"B4",X"09",X"61",X"65",X"67",X"97",X"D0",
		X"0E",X"2A",X"AF",X"C8",X"9A",X"F8",X"18",X"18",X"DB",X"CD",X"CD",X"A0",X"65",X"C7",X"3F",X"21",
		X"71",X"3F",X"65",X"54",X"09",X"65",X"7D",X"3F",X"61",X"2B",X"80",X"38",X"98",X"20",X"99",X"20",
		X"BA",X"A8",X"BB",X"A8",X"A8",X"A8",X"A8",X"A8",X"B8",X"A8",X"B9",X"A8",X"BA",X"A8",X"9B",X"21",
		X"F8",X"EF",X"91",X"51",X"47",X"09",X"07",X"28",X"9E",X"28",X"6D",X"B8",X"61",X"89",X"80",X"29",
		X"AA",X"00",X"88",X"87",X"BA",X"02",X"88",X"26",X"28",X"45",X"BB",X"18",X"A9",X"0C",X"29",X"AA",
		X"80",X"88",X"1E",X"38",X"9A",X"2A",X"20",X"6D",X"13",X"B8",X"61",X"8E",X"90",X"4D",X"8E",X"28",
		X"E1",X"45",X"68",X"2B",X"B2",X"02",X"88",X"DD",X"B6",X"10",X"BA",X"02",X"88",X"45",X"E7",X"2C",
		X"F9",X"92",X"82",X"88",X"65",X"28",X"09",X"B6",X"80",X"6D",X"1C",X"A1",X"65",X"B4",X"09",X"B4",
		X"45",X"3C",X"A1",X"45",X"B4",X"29",X"B4",X"45",X"B4",X"29",X"45",X"3C",X"A1",X"B4",X"45",X"3C",
		X"09",X"6D",X"1C",X"A1",X"65",X"60",X"10",X"49",X"89",X"2A",X"20",X"94",X"04",X"98",X"3E",X"69",
		X"4D",X"2E",X"AB",X"4B",X"AB",X"29",X"B2",X"C0",X"18",X"A7",X"CE",X"0F",X"A0",X"F8",X"41",X"FF",
		X"58",X"07",X"08",X"2E",X"1A",X"B9",X"20",X"07",X"9F",X"68",X"5E",X"83",X"AF",X"A0",X"83",X"F6",
		X"90",X"50",X"F0",X"FF",X"A3",X"BE",X"29",X"87",X"41",X"DB",X"A9",X"60",X"8C",X"2C",X"A0",X"14",
		X"85",X"6D",X"D8",X"B8",X"18",X"AC",X"89",X"71",X"24",X"6D",X"A2",X"B8",X"89",X"09",X"24",X"6D",
		X"0A",X"18",X"D3",X"41",X"BE",X"00",X"87",X"BA",X"70",X"8C",X"BA",X"80",X"8C",X"30",X"53",X"DB",
		X"89",X"18",X"24",X"8C",X"08",X"AD",X"85",X"6D",X"D8",X"B8",X"18",X"2D",X"1E",X"D7",X"9A",X"94",
		X"8C",X"D3",X"41",X"BE",X"28",X"30",X"D2",X"DB",X"A9",X"A0",X"8C",X"2C",X"A0",X"1A",X"2D",X"B2",
		X"C0",X"18",X"0F",X"6B",X"47",X"A0",X"85",X"6D",X"5A",X"B8",X"10",X"2B",X"65",X"70",X"10",X"B0",
		X"2D",X"B6",X"D7",X"BA",X"95",X"8C",X"D3",X"41",X"BE",X"00",X"30",X"FA",X"B6",X"01",X"BA",X"41",
		X"B0",X"69",X"1E",X"28",X"9A",X"69",X"B0",X"69",X"D7",X"46",X"D8",X"FF",X"07",X"0B",X"57",X"F2",
		X"EE",X"27",X"2F",X"83",X"1E",X"28",X"57",X"21",X"3A",X"31",X"11",X"5E",X"8B",X"56",X"65",X"5A",
		X"11",X"61",X"C1",X"28",X"C5",X"28",X"41",X"28",X"45",X"28",X"D2",X"28",X"D7",X"28",X"54",X"28",
		X"EA",X"28",X"EF",X"28",X"E6",X"28",X"FC",X"28",X"F3",X"28",X"0A",X"28",X"02",X"28",X"1A",X"28",
		X"33",X"28",X"AC",X"28",X"2E",X"28",X"39",X"28",X"E4",X"28",X"67",X"28",X"74",X"28",X"69",X"28",
		X"DE",X"28",X"2D",X"29",X"3D",X"29",X"AD",X"29",X"BF",X"29",X"61",X"29",X"75",X"29",X"FA",X"29",
		X"20",X"29",X"37",X"29",X"38",X"29",X"F2",X"29",X"6D",X"29",X"03",X"2A",X"0A",X"2A",X"43",X"2A",
		X"E6",X"2A",X"1B",X"2A",X"92",X"2A",X"CB",X"2A",X"27",X"2B",X"B6",X"2B",X"F8",X"2B",X"8C",X"2B",
		X"73",X"2B",X"96",X"2C",X"D4",X"2C",X"B6",X"2C",X"74",X"2C",X"8E",X"2D",X"DC",X"2D",X"E2",X"2D",
		X"37",X"2E",X"F5",X"2E",X"C8",X"2E",X"60",X"2F",X"9F",X"2F",X"A5",X"20",X"81",X"20",X"A5",X"21",
		X"39",X"A9",X"45",X"AA",X"69",X"AA",X"27",X"AB",X"1F",X"AC",X"7A",X"AC",X"E0",X"AD",X"B1",X"AE",
		X"E7",X"27",X"72",X"38",X"7A",X"39",X"72",X"3A",X"FA",X"3B",X"12",X"3C",X"5B",X"3D",X"37",X"3F",
		X"5F",X"B8",X"FC",X"B9",X"A0",X"BB",X"8A",X"BD",X"76",X"BE",X"BC",X"20",X"AD",X"22",X"BD",X"24",
		X"CC",X"AE",X"BC",X"A1",X"29",X"28",X"29",X"28",X"29",X"28",X"29",X"28",X"29",X"28",X"29",X"28",
		X"81",X"28",X"F5",X"92",X"3E",X"8C",X"91",X"DC",X"11",X"6B",X"27",X"A5",X"EE",X"B9",X"7C",X"B9",
		X"29",X"32",X"2E",X"32",X"23",X"32",X"89",X"29",X"07",X"D1",X"D3",X"77",X"8B",X"0F",X"07",X"0F",
		X"07",X"DF",X"8B",X"D2",X"DF",X"8B",X"07",X"07",X"07",X"07",X"DF",X"61",X"89",X"20",X"27",X"10",
		X"C0",X"A9",X"30",X"8F",X"30",X"E3",X"A9",X"28",X"8F",X"30",X"DE",X"A9",X"B0",X"8F",X"30",X"D9",
		X"63",X"47",X"10",X"2A",X"63",X"67",X"FD",X"B2",X"3E",X"8C",X"91",X"20",X"12",X"4B",X"27",X"A5",
		X"A2",X"1A",X"7B",X"1A",X"F8",X"1A",X"FD",X"1A",X"62",X"1A",X"A9",X"05",X"8F",X"D9",X"43",X"EF",
		X"88",X"A8",X"63",X"E7",X"88",X"39",X"EE",X"AF",X"DF",X"69",X"EE",X"AF",X"C7",X"F6",X"A0",X"76",
		X"AF",X"B0",X"2A",X"B6",X"AF",X"FF",X"41",X"CE",X"AF",X"6F",X"F6",X"18",X"D6",X"0F",X"B0",X"01",
		X"2F",X"D7",X"61",X"81",X"8C",X"8F",X"10",X"5D",X"89",X"34",X"27",X"B8",X"F0",X"81",X"0C",X"8F",
		X"30",X"CB",X"A9",X"3C",X"8F",X"30",X"4E",X"DD",X"B2",X"BE",X"8C",X"39",X"71",X"1A",X"4B",X"8F",
		X"0D",X"F3",X"12",X"0D",X"12",X"8A",X"12",X"8F",X"12",X"1C",X"12",X"81",X"90",X"8F",X"F9",X"46",
		X"2F",X"FF",X"43",X"D6",X"41",X"A9",X"25",X"8F",X"30",X"F4",X"A9",X"35",X"8F",X"30",X"C7",X"A9",
		X"0D",X"8F",X"10",X"C2",X"89",X"B5",X"27",X"B8",X"ED",X"92",X"3E",X"8C",X"75",X"F6",X"80",X"07",
		X"40",X"CE",X"AF",X"D6",X"29",X"44",X"EB",X"1C",X"55",X"BC",X"AB",X"55",X"F6",X"0B",X"55",X"96",
		X"02",X"78",X"75",X"96",X"03",X"28",X"75",X"94",X"01",X"7D",X"63",X"AE",X"C6",X"4C",X"33",X"BC",
		X"55",X"F6",X"A9",X"55",X"96",X"08",X"50",X"55",X"BE",X"09",X"28",X"55",X"F6",X"0C",X"43",X"6F",
		X"08",X"AC",X"75",X"96",X"04",X"28",X"63",X"F7",X"08",X"2C",X"75",X"96",X"06",X"D7",X"75",X"E6",
		X"2A",X"55",X"EE",X"03",X"39",X"E4",X"BA",X"5D",X"F6",X"CD",X"A9",X"2D",X"BB",X"29",X"AB",X"00",
		X"6D",X"11",X"08",X"6C",X"7E",X"D0",X"88",X"B8",X"1E",X"AF",X"75",X"6B",X"06",X"6E",X"08",X"2A",
		X"96",X"D7",X"75",X"77",X"24",X"DD",X"9E",X"26",X"28",X"3E",X"28",X"CD",X"3E",X"32",X"10",X"21",
		X"65",X"D0",X"10",X"75",X"5E",X"AD",X"65",X"3E",X"12",X"E9",X"8B",X"D6",X"75",X"DF",X"00",X"8B",
		X"75",X"75",X"2A",X"DD",X"DC",X"2B",X"79",X"21",X"97",X"04",X"63",X"C6",X"61",X"D7",X"D6",X"D5",
		X"7C",X"D3",X"7A",X"D1",X"FF",X"56",X"FD",X"54",X"63",X"89",X"63",X"18",X"89",X"6D",X"13",X"01",
		X"56",X"23",X"5E",X"EB",X"E1",X"6F",X"34",X"84",X"33",X"B7",X"34",X"BC",X"34",X"A4",X"34",X"73",
		X"13",X"98",X"13",X"02",X"13",X"97",X"13",X"3D",X"14",X"22",X"14",X"75",X"9E",X"28",X"80",X"96",
		X"28",X"CD",X"3E",X"32",X"75",X"36",X"26",X"28",X"89",X"97",X"04",X"CB",X"6E",X"3A",X"96",X"04",
		X"7E",X"2B",X"08",X"2F",X"7E",X"2C",X"08",X"3B",X"E9",X"E9",X"61",X"92",X"91",X"8F",X"FE",X"50",
		X"9A",X"39",X"07",X"21",X"94",X"04",X"9E",X"28",X"E9",X"E1",X"61",X"3A",X"3A",X"07",X"FE",X"D8",
		X"9A",X"3A",X"27",X"89",X"3D",X"8C",X"10",X"C6",X"E9",X"8B",X"5E",X"8B",X"ED",X"65",X"90",X"BA",
		X"E9",X"C9",X"E9",X"23",X"D6",X"23",X"ED",X"CD",X"3C",X"32",X"E9",X"C9",X"E9",X"23",X"75",X"CB",
		X"87",X"F6",X"64",X"C6",X"13",X"65",X"78",X"BB",X"1A",X"93",X"24",X"75",X"DF",X"AA",X"61",X"E9",
		X"8B",X"DD",X"63",X"2E",X"F6",X"CC",X"44",X"33",X"65",X"5E",X"33",X"C9",X"D6",X"DD",X"DF",X"2E",
		X"1D",X"75",X"63",X"2E",X"7E",X"61",X"6B",X"75",X"4E",X"2C",X"75",X"CE",X"85",X"75",X"5E",X"2E",
		X"95",X"DD",X"DF",X"2E",X"EE",X"F7",X"68",X"DD",X"63",X"2E",X"96",X"EB",X"8B",X"C9",X"D6",X"DD",
		X"DF",X"2F",X"1D",X"75",X"63",X"2F",X"7E",X"61",X"ED",X"65",X"48",X"BC",X"E9",X"E3",X"75",X"C6",
		X"2C",X"55",X"EE",X"05",X"55",X"F6",X"2F",X"B5",X"55",X"FF",X"2F",X"CE",X"F7",X"48",X"55",X"43",
		X"87",X"96",X"6B",X"83",X"61",X"41",X"8B",X"F6",X"75",X"D7",X"05",X"83",X"ED",X"6D",X"96",X"BA",
		X"C9",X"41",X"C9",X"AB",X"F6",X"AB",X"CD",X"45",X"67",X"1A",X"C9",X"41",X"C9",X"AB",X"F6",X"AB",
		X"75",X"D7",X"02",X"69",X"E9",X"83",X"5E",X"83",X"75",X"D5",X"84",X"7D",X"DC",X"2D",X"61",X"41",
		X"AB",X"F6",X"AB",X"55",X"FF",X"0E",X"41",X"C9",X"AB",X"AB",X"41",X"45",X"E0",X"1C",X"55",X"FB",
		X"82",X"7D",X"DA",X"2B",X"1A",X"93",X"24",X"7D",X"DF",X"AA",X"75",X"D7",X"03",X"27",X"75",X"D7",
		X"A8",X"55",X"FF",X"06",X"55",X"FF",X"2F",X"41",X"B2",X"BE",X"8C",X"0F",X"3E",X"00",X"77",X"A9",
		X"B1",X"BC",X"11",X"FE",X"8B",X"DE",X"6B",X"7D",X"5E",X"28",X"FE",X"AF",X"75",X"D7",X"80",X"7D",
		X"F6",X"01",X"0F",X"3E",X"28",X"77",X"31",X"76",X"AB",X"7E",X"55",X"FB",X"2C",X"55",X"FA",X"05",
		X"61",X"28",X"D8",X"20",X"D8",X"68",X"D8",X"60",X"D8",X"70",X"D8",X"7D",X"5E",X"A8",X"89",X"13",
		X"BC",X"29",X"A8",X"00",X"C5",X"99",X"43",X"A9",X"43",X"38",X"A9",X"BB",X"BC",X"21",X"76",X"AB",
		X"D6",X"63",X"69",X"38",X"00",X"2C",X"82",X"29",X"10",X"AC",X"86",X"3D",X"15",X"28",X"15",X"C3",
		X"BC",X"CB",X"BC",X"CB",X"BC",X"D0",X"BC",X"D2",X"BC",X"DA",X"BC",X"45",X"40",X"1C",X"30",X"10",
		X"10",X"AE",X"75",X"F6",X"01",X"46",X"81",X"48",X"10",X"2E",X"75",X"F6",X"01",X"46",X"83",X"48",
		X"B6",X"01",X"45",X"14",X"BA",X"A9",X"97",X"8C",X"43",X"4E",X"41",X"55",X"F6",X"09",X"A9",X"E0",
		X"14",X"45",X"7E",X"2D",X"60",X"76",X"02",X"68",X"7E",X"AF",X"60",X"76",X"94",X"68",X"E9",X"69",
		X"75",X"7E",X"21",X"21",X"C8",X"34",X"ED",X"FE",X"2B",X"C8",X"F6",X"2E",X"60",X"FE",X"21",X"C8",
		X"7E",X"AB",X"60",X"E9",X"61",X"75",X"5E",X"A9",X"89",X"40",X"14",X"ED",X"7E",X"2A",X"60",X"F6",
		X"2C",X"C8",X"F6",X"2D",X"60",X"E1",X"61",X"D7",X"D7",X"06",X"2F",X"CD",X"01",X"30",X"96",X"68",
		X"65",X"59",X"08",X"65",X"C8",X"BD",X"65",X"75",X"00",X"0E",X"80",X"18",X"7E",X"65",X"AA",X"BD",
		X"65",X"80",X"35",X"CD",X"86",X"35",X"65",X"9C",X"35",X"CD",X"92",X"35",X"65",X"48",X"35",X"DD",
		X"89",X"00",X"25",X"96",X"85",X"75",X"3E",X"BF",X"88",X"DC",X"1E",X"68",X"65",X"59",X"08",X"61",
		X"75",X"21",X"28",X"05",X"19",X"A8",X"28",X"DD",X"9E",X"37",X"28",X"DD",X"9E",X"2D",X"29",X"DD",
		X"11",X"75",X"9E",X"BF",X"80",X"75",X"9E",X"2D",X"82",X"75",X"11",X"75",X"9E",X"BF",X"80",X"75",
		X"9E",X"2D",X"2B",X"DD",X"11",X"DD",X"9E",X"37",X"28",X"DD",X"9E",X"2D",X"2C",X"DD",X"11",X"DD",
		X"9E",X"BF",X"80",X"75",X"9E",X"2D",X"85",X"75",X"11",X"75",X"9E",X"BF",X"80",X"75",X"9E",X"2D",
		X"2E",X"C9",X"75",X"21",X"28",X"05",X"10",X"34",X"75",X"21",X"A8",X"05",X"10",X"3E",X"75",X"21",
		X"C0",X"8D",X"10",X"38",X"75",X"89",X"C8",X"8D",X"10",X"AA",X"75",X"89",X"A0",X"8D",X"10",X"2C",
		X"75",X"21",X"88",X"05",X"19",X"D1",X"35",X"3A",X"31",X"00",X"AF",X"28",X"25",X"CD",X"07",X"A0",
		X"91",X"41",X"15",X"F6",X"02",X"90",X"83",X"19",X"6D",X"BD",X"75",X"D6",X"17",X"6B",X"27",X"A5",
		X"61",X"2D",X"36",X"C8",X"35",X"4C",X"36",X"54",X"A8",X"4C",X"36",X"C8",X"35",X"7C",X"36",X"C8",
		X"15",X"7A",X"17",X"40",X"15",X"DC",X"88",X"40",X"15",X"9C",X"16",X"40",X"15",X"18",X"17",X"EE",
		X"20",X"E0",X"BD",X"E0",X"BD",X"55",X"BE",X"00",X"28",X"55",X"BE",X"01",X"98",X"55",X"BE",X"02",
		X"00",X"7D",X"5E",X"2D",X"1C",X"B4",X"75",X"D7",X"83",X"6D",X"8E",X"BE",X"75",X"F6",X"85",X"76",
		X"29",X"48",X"55",X"BC",X"BF",X"41",X"55",X"BE",X"2C",X"03",X"55",X"BE",X"2E",X"0A",X"55",X"BE",
		X"87",X"28",X"75",X"96",X"00",X"D7",X"75",X"96",X"01",X"28",X"75",X"96",X"02",X"28",X"75",X"96",
		X"AB",X"00",X"45",X"8F",X"A0",X"27",X"B5",X"55",X"FF",X"1E",X"45",X"AB",X"B1",X"45",X"CE",X"33",
		X"75",X"94",X"17",X"69",X"89",X"0C",X"16",X"6D",X"CC",X"BE",X"75",X"F6",X"85",X"76",X"81",X"48",
		X"55",X"BC",X"BF",X"41",X"55",X"F6",X"2D",X"B5",X"2F",X"2F",X"3E",X"00",X"77",X"31",X"F6",X"AB",
		X"75",X"D7",X"80",X"F6",X"8B",X"7D",X"DF",X"29",X"5E",X"83",X"75",X"D7",X"82",X"F6",X"8B",X"7D",
		X"FF",X"03",X"30",X"A2",X"28",X"98",X"A8",X"09",X"70",X"88",X"70",X"10",X"08",X"88",X"70",X"10",
		X"D8",X"98",X"D8",X"38",X"A0",X"98",X"D8",X"38",X"D8",X"18",X"F8",X"AB",X"89",X"84",X"16",X"6D",
		X"64",X"1E",X"55",X"F6",X"2D",X"D6",X"2C",X"58",X"55",X"BC",X"BF",X"41",X"28",X"28",X"A8",X"0A",
		X"80",X"78",X"00",X"AB",X"80",X"70",X"00",X"29",X"80",X"A8",X"00",X"AB",X"80",X"B8",X"00",X"AD",
		X"28",X"38",X"A8",X"0C",X"45",X"F0",X"BE",X"55",X"BC",X"07",X"55",X"F6",X"2F",X"55",X"96",X"06",
		X"70",X"7D",X"9E",X"2F",X"80",X"B6",X"10",X"7D",X"3E",X"28",X"64",X"3F",X"17",X"B6",X"B8",X"7D",
		X"96",X"00",X"44",X"24",X"BF",X"B6",X"50",X"55",X"96",X"00",X"44",X"4E",X"BF",X"4B",X"5F",X"3D",
		X"1A",X"24",X"20",X"46",X"17",X"48",X"86",X"28",X"75",X"F6",X"17",X"76",X"84",X"80",X"01",X"7D",
		X"D6",X"36",X"F6",X"2B",X"88",X"2A",X"0E",X"B2",X"75",X"34",X"24",X"DD",X"D6",X"24",X"EE",X"2B",
		X"E0",X"75",X"9C",X"AC",X"E3",X"0D",X"19",X"75",X"ED",X"19",X"88",X"28",X"75",X"11",X"75",X"9C",
		X"37",X"DD",X"E9",X"C9",X"75",X"7E",X"2D",X"FE",X"29",X"C0",X"75",X"E5",X"75",X"34",X"37",X"11",
		X"88",X"28",X"75",X"11",X"75",X"9C",X"17",X"75",X"11",X"75",X"9C",X"BF",X"75",X"11",X"75",X"9C",
		X"37",X"DD",X"11",X"DD",X"9C",X"37",X"75",X"19",X"75",X"34",X"37",X"DD",X"E9",X"C9",X"75",X"34",
		X"17",X"61",X"75",X"D6",X"85",X"F6",X"81",X"64",X"F8",X"BE",X"75",X"9C",X"87",X"75",X"5E",X"2F",
		X"75",X"BE",X"2E",X"D8",X"75",X"36",X"2F",X"28",X"96",X"E8",X"75",X"BE",X"28",X"CC",X"F3",X"37",
		X"1E",X"50",X"75",X"B6",X"80",X"64",X"46",X"BF",X"E3",X"5F",X"1D",X"65",X"8C",X"BF",X"75",X"ED",
		X"75",X"21",X"88",X"05",X"75",X"34",X"37",X"DD",X"9C",X"37",X"75",X"E1",X"75",X"35",X"37",X"C9",
		X"65",X"44",X"17",X"75",X"9C",X"2F",X"75",X"D6",X"87",X"75",X"3E",X"2E",X"70",X"75",X"9E",X"2F",
		X"28",X"CD",X"4D",X"37",X"96",X"D7",X"75",X"BE",X"28",X"CC",X"22",X"A8",X"96",X"60",X"75",X"BE",
		X"80",X"64",X"9A",X"20",X"89",X"57",X"17",X"75",X"5E",X"28",X"81",X"3B",X"80",X"E5",X"B9",X"64",
		X"B5",X"A8",X"6B",X"5F",X"B5",X"DD",X"D6",X"2D",X"F6",X"29",X"68",X"DD",X"D6",X"28",X"EE",X"2F",
		X"E0",X"0E",X"96",X"06",X"87",X"75",X"63",X"28",X"56",X"80",X"85",X"65",X"E2",X"EB",X"10",X"2B",
		X"65",X"50",X"63",X"C9",X"75",X"7E",X"2D",X"FE",X"2A",X"CA",X"D8",X"36",X"92",X"AC",X"00",X"E6",
		X"17",X"68",X"86",X"3A",X"E3",X"A8",X"17",X"B0",X"C0",X"E8",X"D0",X"F8",X"C8",X"E0",X"D8",X"F0",
		X"A8",X"28",X"B8",X"38",X"88",X"20",X"98",X"30",X"E8",X"68",X"7D",X"CD",X"7D",X"94",X"37",X"7D",
		X"21",X"C0",X"8D",X"91",X"20",X"88",X"DD",X"9C",X"BF",X"75",X"34",X"BF",X"DD",X"11",X"DD",X"9C",
		X"37",X"7D",X"94",X"BF",X"7D",X"31",X"7D",X"94",X"37",X"7D",X"94",X"BF",X"7D",X"C9",X"6D",X"9D",
		X"2E",X"61",X"DD",X"5E",X"2D",X"7E",X"29",X"60",X"D6",X"8C",X"58",X"E9",X"C9",X"07",X"AF",X"07",
		X"46",X"BF",X"5E",X"8A",X"E7",X"86",X"A6",X"82",X"A0",X"28",X"6D",X"88",X"01",X"69",X"6D",X"44",
		X"BF",X"75",X"34",X"8F",X"DD",X"5E",X"2F",X"75",X"96",X"8E",X"D8",X"75",X"36",X"8F",X"28",X"65",
		X"ED",X"BF",X"7D",X"56",X"A0",X"CE",X"A7",X"6C",X"8C",X"80",X"7D",X"56",X"A0",X"5E",X"41",X"6C",
		X"0D",X"80",X"DD",X"5E",X"28",X"7E",X"A0",X"64",X"1B",X"80",X"DD",X"5E",X"28",X"7E",X"D0",X"64",
		X"38",X"80",X"4B",X"5F",X"15",X"7D",X"F6",X"A9",X"07",X"E8",X"7D",X"96",X"A4",X"8A",X"7D",X"96",
		X"A9",X"77",X"C9",X"75",X"36",X"8C",X"2B",X"61",X"DD",X"9C",X"BF",X"75",X"F6",X"8D",X"D6",X"8E",
		X"7D",X"94",X"37",X"69",X"7D",X"56",X"A0",X"27",X"AF",X"27",X"46",X"BF",X"5E",X"89",X"76",X"8B",
		X"D8",X"7E",X"B8",X"F0",X"E7",X"8E",X"29",X"8A",X"28",X"28",X"B6",X"AE",X"DD",X"63",X"2C",X"CE",
		X"80",X"8A",X"B6",X"88",X"8E",X"A8",X"4D",X"6D",X"05",X"A1",X"6D",X"B9",X"01",X"E9",X"98",X"56",
		X"C9",X"8E",X"28",X"75",X"E6",X"BE",X"A1",X"11",X"FE",X"8B",X"7E",X"61",X"39",X"60",X"20",X"65",
		X"F9",X"80",X"7D",X"56",X"23",X"EB",X"2F",X"A5",X"58",X"80",X"64",X"81",X"A8",X"81",X"18",X"81",
		X"CC",X"81",X"65",X"82",X"CC",X"81",X"65",X"82",X"30",X"81",X"D2",X"B7",X"E6",X"C8",X"BF",X"C8",
		X"46",X"48",X"5A",X"97",X"46",X"48",X"37",X"48",X"46",X"48",X"10",X"89",X"5A",X"97",X"46",X"48",
		X"BF",X"40",X"E6",X"40",X"D2",X"3F",X"E6",X"40",X"BF",X"40",X"E6",X"40",X"68",X"21",X"D2",X"3F",
		X"46",X"48",X"37",X"48",X"46",X"48",X"5A",X"97",X"46",X"48",X"37",X"48",X"46",X"48",X"60",X"89",
		X"DD",X"36",X"2C",X"01",X"DD",X"34",X"AB",X"C9",X"DD",X"36",X"2C",X"02",X"DD",X"34",X"AB",X"C9",
		X"75",X"36",X"A4",X"0B",X"75",X"34",X"23",X"C9",X"75",X"34",X"37",X"C9",X"E0",X"89",X"5A",X"97",
		X"E6",X"40",X"BF",X"40",X"E6",X"40",X"D2",X"3F",X"E6",X"40",X"BF",X"40",X"E6",X"40",X"70",X"21",
		X"46",X"48",X"54",X"89",X"46",X"48",X"D0",X"89",X"46",X"48",X"54",X"89",X"46",X"48",X"60",X"89",
		X"2E",X"78",X"DD",X"70",X"2A",X"CD",X"83",X"39",X"DD",X"34",X"AB",X"C9",X"2E",X"7C",X"B8",X"F2",
		X"2E",X"89",X"8A",X"89",X"2E",X"89",X"0D",X"89",X"2E",X"89",X"E0",X"89",X"60",X"89",X"75",X"CB",
		X"A9",X"46",X"CC",X"99",X"21",X"CD",X"0A",X"40",X"C9",X"DD",X"36",X"0A",X"AA",X"DD",X"36",X"09",
		X"27",X"C9",X"75",X"36",X"A2",X"3C",X"65",X"A3",X"11",X"DD",X"9C",X"03",X"61",X"DD",X"9E",X"0A",
		X"3A",X"CD",X"83",X"39",X"DD",X"34",X"AB",X"C9",X"8E",X"21",X"30",X"21",X"8E",X"21",X"68",X"21",
		X"EC",X"89",X"60",X"89",X"75",X"36",X"24",X"08",X"75",X"34",X"23",X"C9",X"E0",X"8A",X"2E",X"89",
		X"AC",X"22",X"E6",X"40",X"BB",X"22",X"E6",X"40",X"AC",X"22",X"E6",X"40",X"BB",X"22",X"8E",X"21",
		X"24",X"8A",X"46",X"48",X"33",X"8A",X"46",X"48",X"24",X"8A",X"46",X"48",X"33",X"8A",X"2E",X"89",
		X"8E",X"21",X"A2",X"22",X"8E",X"21",X"35",X"22",X"AC",X"22",X"E6",X"40",X"BB",X"22",X"E6",X"40",
		X"24",X"82",X"46",X"C8",X"33",X"82",X"2E",X"81",X"BF",X"82",X"60",X"81",X"7D",X"96",X"A0",X"D2",
		X"DD",X"9E",X"29",X"1A",X"CD",X"6E",X"33",X"75",X"34",X"AB",X"C9",X"75",X"36",X"88",X"70",X"75",
		X"96",X"89",X"B8",X"6D",X"6E",X"93",X"7D",X"94",X"23",X"69",X"7D",X"96",X"A2",X"54",X"6D",X"23",
		X"B1",X"75",X"34",X"AB",X"C9",X"75",X"36",X"8A",X"50",X"65",X"83",X"B1",X"DD",X"9C",X"AB",X"61",
		X"86",X"9B",X"A6",X"AC",X"82",X"88",X"28",X"16",X"B2",X"92",X"A2",X"28",X"B6",X"18",X"8E",X"8C",
		X"CD",X"B4",X"A1",X"1C",X"38",X"72",X"CD",X"83",X"A1",X"86",X"2C",X"65",X"B4",X"A1",X"B4",X"90",
		X"5A",X"7D",X"94",X"AB",X"69",X"C8",X"82",X"1F",X"82",X"2E",X"81",X"2E",X"81",X"2E",X"81",X"06",
		X"22",X"15",X"22",X"E6",X"68",X"48",X"22",X"E6",X"68",X"15",X"22",X"E6",X"68",X"1F",X"22",X"2E",
		X"81",X"2E",X"81",X"06",X"82",X"15",X"82",X"E6",X"E0",X"48",X"82",X"2E",X"81",X"2E",X"81",X"15",
		X"22",X"E6",X"68",X"1F",X"22",X"E8",X"21",X"75",X"36",X"88",X"28",X"75",X"36",X"89",X"28",X"65",
		X"6E",X"93",X"7D",X"94",X"23",X"69",X"7D",X"96",X"A0",X"F6",X"7D",X"96",X"A1",X"28",X"6D",X"6E",
		X"33",X"75",X"34",X"AB",X"C9",X"75",X"36",X"8A",X"C0",X"65",X"83",X"B1",X"DD",X"9C",X"AB",X"61",
		X"7D",X"96",X"A2",X"64",X"6D",X"23",X"11",X"7D",X"94",X"AB",X"69",X"6D",X"31",X"83",X"6D",X"85",
		X"23",X"65",X"60",X"BD",X"CD",X"D5",X"A8",X"86",X"28",X"90",X"D6",X"90",X"D6",X"1A",X"24",X"28",
		X"07",X"80",X"A6",X"12",X"85",X"28",X"6D",X"74",X"84",X"6D",X"16",X"83",X"6D",X"CC",X"83",X"6D",
		X"EA",X"83",X"CD",X"D8",X"23",X"65",X"7E",X"83",X"CD",X"FC",X"23",X"75",X"F6",X"BF",X"D6",X"8A",
		X"88",X"7A",X"96",X"48",X"65",X"79",X"00",X"CD",X"4C",X"8C",X"65",X"06",X"83",X"C9",X"A7",X"32",
		X"6F",X"90",X"32",X"42",X"18",X"32",X"6E",X"90",X"C9",X"B6",X"29",X"32",X"6F",X"90",X"32",X"42",
		X"B8",X"32",X"E6",X"38",X"61",X"21",X"A0",X"2C",X"19",X"09",X"AC",X"29",X"5E",X"0B",X"9E",X"18",
		X"C5",X"10",X"21",X"00",X"60",X"39",X"28",X"80",X"29",X"00",X"2C",X"C5",X"10",X"C9",X"DD",X"21",
		X"A0",X"25",X"10",X"14",X"75",X"21",X"80",X"25",X"10",X"1E",X"75",X"21",X"E0",X"25",X"10",X"18",
		X"DD",X"21",X"60",X"8D",X"B8",X"0A",X"DD",X"21",X"08",X"8D",X"B8",X"04",X"DD",X"21",X"00",X"8D",
		X"75",X"F6",X"37",X"39",X"41",X"8B",X"6B",X"27",X"05",X"DB",X"83",X"EF",X"83",X"C7",X"83",X"CD",
		X"D7",X"23",X"C9",X"21",X"17",X"23",X"DD",X"F6",X"2D",X"B5",X"0F",X"0F",X"0F",X"3E",X"28",X"FF",
		X"11",X"F6",X"75",X"77",X"A0",X"23",X"D6",X"DD",X"DF",X"09",X"8B",X"F6",X"2F",X"0F",X"75",X"77",
		X"2A",X"23",X"F6",X"DD",X"77",X"03",X"23",X"F6",X"DD",X"77",X"2C",X"23",X"F6",X"DD",X"77",X"06",
		X"8B",X"DD",X"9E",X"0F",X"A0",X"F6",X"75",X"77",X"B0",X"23",X"D6",X"DD",X"DF",X"19",X"8B",X"DD",
		X"36",X"12",X"28",X"DD",X"34",X"1F",X"C9",X"78",X"78",X"0E",X"2A",X"01",X"AC",X"00",X"E0",X"78",
		X"F0",X"06",X"A3",X"09",X"24",X"08",X"43",X"D0",X"F0",X"06",X"A4",X"09",X"24",X"08",X"41",X"D0",
		X"78",X"0E",X"2D",X"01",X"AC",X"20",X"E2",X"78",X"78",X"0E",X"A8",X"01",X"AC",X"00",X"E5",X"78",
		X"F0",X"06",X"24",X"09",X"24",X"08",X"46",X"CD",X"5F",X"8B",X"75",X"34",X"A7",X"DD",X"D6",X"0F",
		X"DD",X"96",X"2E",X"D8",X"DD",X"36",X"2F",X"00",X"CD",X"35",X"24",X"CD",X"00",X"24",X"C9",X"B2",
		X"84",X"28",X"46",X"8F",X"48",X"7D",X"94",X"AC",X"7D",X"56",X"A2",X"CE",X"58",X"7D",X"6B",X"AC",
		X"7E",X"88",X"2A",X"63",X"5F",X"75",X"77",X"8A",X"DD",X"5E",X"2C",X"7E",X"2B",X"88",X"2C",X"75",
		X"6B",X"8A",X"6E",X"7D",X"6B",X"9A",X"E6",X"00",X"A4",X"7D",X"6B",X"8A",X"6E",X"6D",X"0B",X"B1",
		X"C9",X"65",X"0D",X"B1",X"C9",X"75",X"E6",X"98",X"DD",X"CE",X"39",X"5E",X"6F",X"EE",X"48",X"88",
		X"26",X"50",X"46",X"8F",X"7D",X"D7",X"A4",X"83",X"7D",X"D5",X"B0",X"7D",X"D4",X"99",X"69",X"A7",
		X"2F",X"EE",X"2B",X"91",X"E0",X"84",X"CD",X"2F",X"A5",X"75",X"E6",X"98",X"DD",X"CE",X"39",X"8B",
		X"7D",X"D5",X"B0",X"7D",X"D4",X"99",X"B8",X"6D",X"3F",X"84",X"D5",X"84",X"2E",X"84",X"D0",X"84",
		X"DD",X"9C",X"BF",X"E9",X"C9",X"75",X"E6",X"98",X"DD",X"CE",X"39",X"5E",X"0F",X"A7",X"0F",X"75",
		X"D7",X"8A",X"7D",X"96",X"B2",X"88",X"6B",X"46",X"68",X"7D",X"96",X"9A",X"5F",X"69",X"7D",X"46",
		X"38",X"75",X"66",X"99",X"F6",X"EE",X"AF",X"75",X"77",X"8E",X"DD",X"9E",X"2F",X"88",X"C9",X"61",
		X"81",X"35",X"84",X"CD",X"7D",X"56",X"A4",X"B1",X"0D",X"84",X"4B",X"2F",X"05",X"48",X"84",X"4C",
		X"24",X"68",X"24",X"6C",X"24",X"58",X"24",X"5F",X"24",X"7E",X"24",X"45",X"24",X"E3",X"CE",X"93",
		X"7D",X"95",X"A1",X"69",X"7D",X"94",X"A1",X"69",X"7D",X"95",X"A0",X"69",X"7D",X"94",X"A0",X"69",
		X"CD",X"48",X"24",X"65",X"CC",X"84",X"C9",X"65",X"48",X"84",X"CD",X"68",X"24",X"61",X"CD",X"4C",
		X"84",X"6D",X"6C",X"84",X"69",X"6D",X"EC",X"84",X"6D",X"68",X"84",X"69",X"8E",X"AC",X"4D",X"50",
		X"CD",X"74",X"24",X"1E",X"A9",X"65",X"59",X"A0",X"49",X"90",X"53",X"61",X"46",X"AF",X"56",X"98",
		X"89",X"48",X"AC",X"39",X"B5",X"08",X"06",X"14",X"0E",X"03",X"DF",X"23",X"18",X"F4",X"11",X"AD",
		X"20",X"F6",X"21",X"C0",X"0F",X"2E",X"B7",X"77",X"23",X"38",X"D4",X"C9",X"7B",X"4E",X"EF",X"2D",
		X"E2",X"4D",X"E5",X"88",X"E4",X"41",X"F3",X"58",X"64",X"49",X"71",X"88",X"80",X"4A",X"71",X"88",
		X"EE",X"41",X"EB",X"41",X"EB",X"55",X"ED",X"41",X"20",X"41",X"EB",X"49",X"7A",X"41",X"D7",X"FF",
		X"89",X"78",X"A7",X"22",X"70",X"20",X"8A",X"5A",X"28",X"22",X"64",X"20",X"8A",X"4E",X"28",X"22",
		X"68",X"88",X"21",X"42",X"88",X"39",X"2E",X"00",X"B6",X"01",X"2E",X"05",X"77",X"B9",X"38",X"FC",
		X"89",X"53",X"28",X"B6",X"E1",X"CD",X"29",X"8D",X"89",X"5D",X"28",X"B6",X"63",X"CD",X"29",X"8D",
		X"21",X"4F",X"88",X"B6",X"E9",X"CD",X"89",X"25",X"21",X"49",X"88",X"B6",X"7A",X"CD",X"89",X"25",
		X"89",X"4B",X"28",X"B6",X"E1",X"CD",X"29",X"8D",X"61",X"77",X"8B",X"77",X"8B",X"77",X"61",X"CD",
		X"E8",X"26",X"B2",X"5F",X"88",X"D6",X"2E",X"C8",X"CD",X"E5",X"A0",X"CD",X"17",X"31",X"2E",X"09",
		X"65",X"21",X"30",X"CD",X"3E",X"8E",X"89",X"12",X"00",X"2E",X"20",X"CD",X"53",X"8F",X"89",X"0E",
		X"2E",X"22",X"28",X"88",X"B6",X"10",X"32",X"02",X"88",X"CD",X"8D",X"26",X"C3",X"CD",X"68",X"2B",
		X"65",X"5C",X"04",X"B6",X"90",X"CD",X"14",X"81",X"89",X"07",X"A6",X"22",X"A0",X"20",X"65",X"27",
		X"A0",X"26",X"28",X"E7",X"CD",X"40",X"A3",X"CD",X"E7",X"2C",X"21",X"16",X"2E",X"22",X"28",X"88",
		X"96",X"49",X"0E",X"0B",X"65",X"94",X"01",X"38",X"5B",X"B2",X"77",X"20",X"95",X"6F",X"2F",X"08",
		X"4E",X"0E",X"7F",X"BE",X"3E",X"5D",X"D5",X"41",X"DD",X"21",X"3E",X"06",X"BE",X"02",X"C5",X"7B",
		X"A0",X"28",X"B6",X"B8",X"8E",X"9F",X"6D",X"A5",X"01",X"B0",X"5B",X"12",X"77",X"28",X"CF",X"16",
		X"2D",X"B0",X"0F",X"C7",X"0F",X"A0",X"3E",X"88",X"FF",X"89",X"6B",X"28",X"B9",X"ED",X"CD",X"6F",
		X"86",X"C9",X"B2",X"FE",X"28",X"D7",X"83",X"7D",X"83",X"5D",X"83",X"CD",X"6D",X"6F",X"86",X"C9",
		X"B2",X"FE",X"88",X"DF",X"23",X"75",X"23",X"7D",X"23",X"ED",X"CD",X"6F",X"26",X"E9",X"B2",X"FE",
		X"28",X"D7",X"B6",X"08",X"6D",X"59",X"00",X"69",X"B6",X"8E",X"92",X"FF",X"28",X"6D",X"2D",X"86",
		X"A2",X"C8",X"88",X"65",X"99",X"A5",X"58",X"1E",X"2D",X"9A",X"FF",X"28",X"A2",X"CE",X"88",X"65",
		X"39",X"A5",X"58",X"16",X"A4",X"92",X"77",X"28",X"A2",X"EC",X"28",X"6D",X"39",X"A5",X"58",X"16",
		X"2B",X"9A",X"FF",X"28",X"A2",X"DA",X"88",X"65",X"99",X"A5",X"58",X"1E",X"2A",X"9A",X"FF",X"28",
		X"A2",X"F8",X"28",X"6D",X"39",X"A5",X"58",X"16",X"A1",X"92",X"77",X"28",X"69",X"12",X"B6",X"28",
		X"CB",X"C7",X"A0",X"8D",X"C5",X"53",X"38",X"28",X"C9",X"6D",X"FB",X"AE",X"88",X"61",X"39",X"C8",
		X"28",X"81",X"E6",X"28",X"B2",X"FF",X"28",X"E7",X"B6",X"8D",X"18",X"00",X"21",X"AF",X"CF",X"AF",
		X"08",X"86",X"28",X"47",X"C5",X"B8",X"C3",X"ED",X"CD",X"2D",X"26",X"E9",X"73",X"8B",X"72",X"8B",
		X"45",X"6D",X"2F",X"A0",X"41",X"D7",X"83",X"16",X"80",X"D7",X"83",X"D7",X"83",X"D7",X"69",X"16",
		X"38",X"9A",X"2A",X"28",X"21",X"FE",X"88",X"9E",X"69",X"65",X"7E",X"87",X"B6",X"AA",X"CD",X"59",
		X"00",X"A6",X"24",X"ED",X"6D",X"73",X"02",X"07",X"49",X"CE",X"2C",X"00",X"A7",X"16",X"A1",X"6D",
		X"59",X"A0",X"38",X"67",X"CD",X"73",X"A2",X"0F",X"CB",X"5F",X"20",X"EE",X"CB",X"D7",X"20",X"90",
		X"63",X"FF",X"88",X"91",X"92",X"C8",X"2C",X"07",X"88",X"00",X"E9",X"41",X"96",X"48",X"65",X"79",
		X"A0",X"C9",X"CD",X"75",X"A8",X"B2",X"25",X"88",X"46",X"07",X"20",X"D8",X"2E",X"10",X"B2",X"25",
		X"28",X"CB",X"57",X"20",X"A2",X"2E",X"B6",X"F0",X"9A",X"0A",X"28",X"CD",X"F6",X"8F",X"10",X"6C",
		X"21",X"5E",X"88",X"35",X"B6",X"40",X"96",X"20",X"00",X"36",X"FB",X"B8",X"9C",X"21",X"FE",X"88",
		X"9C",X"B6",X"74",X"96",X"88",X"3B",X"9E",X"49",X"10",X"27",X"65",X"CB",X"87",X"B6",X"30",X"32",
		X"2A",X"88",X"CD",X"56",X"27",X"C9",X"DD",X"45",X"41",X"22",X"28",X"88",X"B2",X"5E",X"88",X"CD",
		X"14",X"81",X"61",X"B6",X"30",X"32",X"A2",X"20",X"F5",X"45",X"10",X"E4",X"89",X"FF",X"87",X"2E",
		X"2A",X"CD",X"54",X"29",X"38",X"FB",X"21",X"45",X"A0",X"2E",X"2E",X"CD",X"54",X"29",X"38",X"FB",
		X"96",X"19",X"9A",X"0A",X"28",X"39",X"A6",X"06",X"89",X"50",X"28",X"CD",X"9B",X"8F",X"19",X"0E",
		X"39",X"21",X"7A",X"88",X"CD",X"B3",X"27",X"39",X"2E",X"14",X"21",X"4C",X"88",X"CD",X"13",X"27",
		X"19",X"0E",X"B7",X"21",X"E6",X"20",X"65",X"BB",X"87",X"39",X"A6",X"12",X"89",X"48",X"28",X"CD",
		X"13",X"27",X"C9",X"C5",X"7B",X"00",X"88",X"FE",X"23",X"7E",X"23",X"45",X"C3",X"CD",X"68",X"2B",
		X"65",X"5C",X"04",X"B6",X"90",X"CD",X"14",X"81",X"0E",X"0B",X"65",X"08",X"01",X"38",X"5B",X"41",
		X"F6",X"23",X"45",X"26",X"28",X"E7",X"CD",X"40",X"A3",X"CD",X"E7",X"2C",X"2E",X"05",X"CD",X"00",
		X"01",X"38",X"5B",X"41",X"65",X"E0",X"87",X"C9",X"D6",X"CD",X"14",X"81",X"8B",X"F6",X"65",X"94",
		X"A1",X"23",X"F6",X"CD",X"B4",X"29",X"C9",X"07",X"A8",X"18",X"7C",X"4F",X"6C",X"41",X"F9",X"3E",
		X"F3",X"80",X"80",X"CA",X"E5",X"DB",X"F4",X"80",X"9D",X"8F",X"A5",X"98",X"64",X"E9",X"F3",X"DC",
		X"20",X"EF",X"6E",X"80",X"78",X"EC",X"69",X"F9",X"6D",X"5A",X"2D",X"8A",X"B8",X"CD",X"EE",X"DC",
		X"E5",X"DA",X"80",X"F9",X"67",X"DD",X"F2",X"80",X"61",X"EE",X"61",X"DC",X"61",X"C9",X"64",X"5B",
		X"2F",X"8C",X"3F",X"DB",X"6B",X"EF",X"7A",X"CD",X"20",X"80",X"20",X"C9",X"6B",X"DC",X"20",X"80",
		X"80",X"EE",X"E1",X"ED",X"ED",X"8F",X"23",X"B9",X"F3",X"CB",X"67",X"DA",X"E5",X"80",X"80",X"80",
		X"69",X"CB",X"7C",X"80",X"20",X"80",X"EE",X"C9",X"ED",X"4D",X"2A",X"AE",X"39",X"91",X"7B",X"5C",
		X"A2",X"99",X"B1",X"92",X"66",X"4C",X"A2",X"9C",X"B1",X"93",X"F2",X"4C",X"A2",X"9F",X"B1",X"94",
		X"7C",X"68",X"2A",X"BA",X"39",X"95",X"7C",X"68",X"2E",X"88",X"B2",X"B8",X"88",X"63",X"6F",X"08",
		X"21",X"12",X"B6",X"28",X"6B",X"E7",X"A0",X"8A",X"8E",X"77",X"F0",X"92",X"E3",X"18",X"69",X"81",
		X"3A",X"28",X"B2",X"9E",X"88",X"63",X"6F",X"08",X"2B",X"89",X"3B",X"28",X"F6",X"61",X"21",X"9C",
		X"28",X"12",X"B6",X"28",X"6B",X"E7",X"A0",X"8B",X"81",X"9D",X"28",X"56",X"46",X"F7",X"69",X"12",
		X"B9",X"28",X"07",X"60",X"B2",X"9E",X"88",X"63",X"6F",X"08",X"AB",X"0A",X"38",X"28",X"B9",X"8A",
		X"B0",X"28",X"6D",X"84",X"04",X"69",X"A2",X"AE",X"28",X"31",X"82",X"AE",X"28",X"6D",X"0E",X"A3",
		X"C9",X"9A",X"20",X"28",X"B2",X"80",X"88",X"AF",X"20",X"72",X"C9",X"9A",X"21",X"28",X"B2",X"81",
		X"28",X"8F",X"80",X"72",X"69",X"81",X"A0",X"08",X"99",X"89",X"A8",X"A1",X"5E",X"8B",X"96",X"80",
		X"C5",X"B8",X"21",X"88",X"0C",X"91",X"29",X"0C",X"29",X"76",X"2B",X"9E",X"28",X"6D",X"10",X"61",
		X"FD",X"B6",X"80",X"CD",X"14",X"81",X"F9",X"C9",X"6D",X"2E",X"A3",X"55",X"ED",X"21",X"A0",X"20",
		X"F6",X"18",X"77",X"23",X"34",X"41",X"51",X"49",X"C9",X"4D",X"2E",X"01",X"B8",X"ED",X"4D",X"2E",
		X"A2",X"B8",X"48",X"4D",X"0E",X"0C",X"10",X"EB",X"6D",X"2E",X"32",X"B8",X"7E",X"55",X"6D",X"5D",
		X"45",X"55",X"C5",X"EB",X"28",X"88",X"CD",X"6F",X"A1",X"51",X"B8",X"13",X"55",X"4D",X"5D",X"45",
		X"FD",X"C5",X"43",X"08",X"28",X"CD",X"47",X"81",X"F9",X"77",X"92",X"0A",X"28",X"46",X"37",X"39",
		X"28",X"04",X"B9",X"77",X"F1",X"B4",X"EF",X"D6",X"BD",X"B0",X"AB",X"AE",X"28",X"F0",X"B4",X"6F",
		X"F6",X"8C",X"90",X"0A",X"0E",X"08",X"E5",X"6B",X"A0",X"20",X"E9",X"59",X"69",X"51",X"61",X"F0",
		X"D6",X"20",X"30",X"15",X"F1",X"D6",X"BC",X"30",X"B1",X"0F",X"3E",X"00",X"FF",X"21",X"16",X"29",
		X"11",X"FE",X"8B",X"7E",X"8E",X"08",X"C0",X"B9",X"61",X"D6",X"82",X"30",X"24",X"21",X"A2",X"28",
		X"CB",X"6F",X"A0",X"03",X"21",X"22",X"08",X"B8",X"AE",X"D6",X"24",X"30",X"3D",X"21",X"4A",X"83",
		X"63",X"6F",X"80",X"0B",X"89",X"EA",X"AB",X"B6",X"33",X"91",X"90",X"0E",X"39",X"3E",X"A0",X"FF",
		X"B9",X"C9",X"21",X"00",X"08",X"C9",X"00",X"83",X"08",X"83",X"60",X"83",X"68",X"83",X"20",X"83",
		X"A0",X"2B",X"C8",X"2A",X"E8",X"2A",X"88",X"2A",X"A8",X"2A",X"C0",X"2A",X"E0",X"2A",X"80",X"2A",
		X"28",X"82",X"40",X"81",X"48",X"81",X"00",X"81",X"08",X"81",X"60",X"81",X"68",X"81",X"20",X"81",
		X"A0",X"29",X"C8",X"28",X"E8",X"28",X"88",X"28",X"A8",X"28",X"C0",X"28",X"E0",X"28",X"80",X"28",
		X"28",X"80",X"28",X"80",X"F6",X"32",X"28",X"88",X"23",X"F6",X"32",X"01",X"88",X"23",X"F6",X"32",
		X"A2",X"28",X"83",X"56",X"6B",X"57",X"80",X"9A",X"6D",X"B4",X"01",X"83",X"B2",X"8A",X"28",X"6B",
		X"F7",X"08",X"50",X"1E",X"2C",X"65",X"59",X"A0",X"B8",X"61",X"46",X"F7",X"CD",X"B4",X"A1",X"8B",
		X"B2",X"8A",X"28",X"6B",X"F7",X"68",X"B6",X"8C",X"6D",X"59",X"00",X"69",X"81",X"F5",X"02",X"6D",
		X"54",X"A1",X"21",X"0F",X"A2",X"65",X"54",X"A1",X"29",X"1F",X"A2",X"96",X"29",X"1A",X"A8",X"28",
		X"32",X"80",X"A3",X"A1",X"08",X"A2",X"C0",X"41",X"6D",X"54",X"01",X"81",X"18",X"A2",X"6D",X"54",
		X"A1",X"65",X"F2",X"A3",X"21",X"6E",X"A2",X"65",X"54",X"A1",X"21",X"7C",X"A2",X"65",X"54",X"A1",
		X"81",X"53",X"02",X"12",X"E0",X"18",X"6B",X"E7",X"4C",X"54",X"01",X"16",X"23",X"92",X"A2",X"28",
		X"26",X"9C",X"A6",X"8B",X"22",X"88",X"88",X"1E",X"24",X"65",X"28",X"A7",X"C9",X"AA",X"A9",X"9F",
		X"F0",X"80",X"F5",X"80",X"F3",X"80",X"68",X"8F",X"24",X"98",X"F3",X"DC",X"E1",X"DA",X"F4",X"80",
		X"20",X"CA",X"7D",X"DC",X"7C",X"EF",X"CE",X"8F",X"AF",X"B8",X"31",X"80",X"EF",X"DA",X"20",X"92",
		X"80",X"D8",X"64",X"C9",X"71",X"CD",X"F2",X"5B",X"A7",X"AF",X"30",X"91",X"80",X"D8",X"64",X"C9",
		X"F9",X"CD",X"7A",X"80",X"EF",X"EE",X"EC",X"79",X"2F",X"9A",X"38",X"CB",X"7A",X"CD",X"6C",X"E9",
		X"F4",X"00",X"A7",X"AF",X"B0",X"CE",X"F2",X"CD",X"E5",X"80",X"F0",X"EC",X"E1",X"79",X"20",X"B9",
		X"38",X"C8",X"20",X"DB",X"6D",X"CF",X"69",X"80",X"31",X"B1",X"B0",X"12",X"2E",X"9D",X"B8",X"CA",
		X"67",X"EE",X"F5",X"DB",X"80",X"CE",X"67",X"DA",X"80",X"93",X"90",X"90",X"90",X"90",X"80",X"D8",
		X"7C",X"DB",X"92",X"98",X"3D",X"B8",X"35",X"90",X"30",X"90",X"10",X"1A",X"B8",X"28",X"07",X"08",
		X"23",X"B2",X"B6",X"20",X"EE",X"09",X"80",X"0C",X"92",X"28",X"B8",X"C9",X"92",X"68",X"B8",X"C9",
		X"21",X"20",X"A3",X"CD",X"54",X"29",X"CD",X"93",X"A3",X"CD",X"86",X"2B",X"CD",X"24",X"A4",X"C9",
		X"A1",X"8A",X"B1",X"99",X"F0",X"88",X"80",X"88",X"80",X"88",X"80",X"88",X"60",X"41",X"80",X"88",
		X"20",X"20",X"20",X"20",X"20",X"32",X"58",X"01",X"21",X"10",X"6B",X"52",X"6D",X"44",X"E9",X"D4",
		X"75",X"45",X"F5",X"45",X"F5",X"21",X"D0",X"83",X"75",X"21",X"A3",X"20",X"A7",X"D5",X"56",X"08",
		X"D5",X"7E",X"29",X"07",X"C5",X"7A",X"B0",X"03",X"B4",X"B8",X"D0",X"B9",X"56",X"30",X"DD",X"77",
		X"A0",X"DD",X"8B",X"D5",X"8B",X"D5",X"8B",X"CB",X"4B",X"A0",X"C9",X"D5",X"E9",X"DD",X"E9",X"C9",
		X"38",X"27",X"C0",X"03",X"64",X"00",X"AA",X"00",X"29",X"00",X"B2",X"08",X"88",X"26",X"28",X"E7",
		X"65",X"48",X"03",X"26",X"B2",X"A6",X"27",X"22",X"A0",X"20",X"96",X"18",X"9A",X"0A",X"28",X"CD",
		X"E7",X"2C",X"C9",X"A2",X"AC",X"88",X"CD",X"40",X"A3",X"26",X"22",X"A6",X"AC",X"22",X"28",X"88",
		X"96",X"18",X"9A",X"0A",X"28",X"CD",X"F4",X"84",X"96",X"98",X"65",X"94",X"01",X"C9",X"82",X"06",
		X"88",X"CD",X"68",X"2B",X"26",X"22",X"A6",X"03",X"22",X"00",X"88",X"B6",X"38",X"32",X"2A",X"88",
		X"65",X"5C",X"04",X"B6",X"90",X"CD",X"14",X"81",X"65",X"76",X"03",X"A2",X"24",X"20",X"E5",X"FB",
		X"AE",X"88",X"CD",X"99",X"A5",X"58",X"C5",X"7B",X"AC",X"88",X"CD",X"93",X"A3",X"C9",X"21",X"14",
		X"28",X"CB",X"D6",X"48",X"ED",X"A2",X"26",X"20",X"19",X"B0",X"23",X"B2",X"E0",X"38",X"63",X"6F",
		X"A0",X"03",X"39",X"88",X"3B",X"CD",X"99",X"2D",X"41",X"D8",X"34",X"CB",X"D6",X"CD",X"3B",X"2D",
		X"8E",X"89",X"6D",X"27",X"30",X"69",X"81",X"9D",X"28",X"6B",X"F6",X"E8",X"45",X"02",X"B0",X"28",
		X"39",X"30",X"AB",X"1A",X"68",X"18",X"CB",X"C7",X"A0",X"8B",X"39",X"28",X"3B",X"65",X"99",X"A5",
		X"41",X"78",X"B8",X"5E",X"A2",X"98",X"28",X"6D",X"E0",X"A3",X"86",X"82",X"A6",X"9D",X"82",X"88",
		X"88",X"1E",X"38",X"9A",X"2A",X"28",X"CD",X"DC",X"A4",X"1E",X"30",X"65",X"B4",X"A1",X"CD",X"8E",
		X"04",X"02",X"24",X"28",X"65",X"73",X"B0",X"28",X"6D",X"39",X"05",X"F8",X"65",X"F3",X"24",X"28",
		X"CD",X"1B",X"A3",X"61",X"2E",X"8D",X"21",X"8B",X"88",X"5E",X"D6",X"90",X"20",X"A9",X"B6",X"80",
		X"6D",X"B4",X"01",X"83",X"98",X"53",X"69",X"56",X"6D",X"B4",X"01",X"83",X"98",X"71",X"69",X"A6",
		X"2A",X"89",X"2E",X"28",X"B8",X"43",X"21",X"54",X"A4",X"65",X"54",X"A1",X"21",X"8A",X"A5",X"65",
		X"DC",X"A1",X"6D",X"2F",X"00",X"86",X"A0",X"47",X"6D",X"C8",X"03",X"6D",X"47",X"A4",X"81",X"8F",
		X"21",X"8A",X"28",X"28",X"B6",X"AA",X"32",X"8A",X"88",X"65",X"8F",X"A0",X"D6",X"8E",X"B0",X"8C",
		X"5E",X"8D",X"B8",X"70",X"CF",X"ED",X"B6",X"AE",X"6D",X"B4",X"01",X"16",X"27",X"6D",X"14",X"A1",
		X"49",X"90",X"52",X"86",X"28",X"65",X"8F",X"A0",X"D6",X"8E",X"B0",X"8D",X"5E",X"8D",X"2C",X"10",
		X"DF",X"A5",X"8C",X"68",X"4D",X"50",X"B5",X"B6",X"A0",X"77",X"81",X"A8",X"05",X"31",X"F6",X"86",
		X"23",X"4F",X"22",X"88",X"88",X"ED",X"B6",X"A8",X"CD",X"B4",X"A1",X"1E",X"A9",X"65",X"B4",X"A1",
		X"41",X"86",X"A0",X"82",X"A0",X"28",X"B6",X"AA",X"6D",X"B4",X"01",X"16",X"23",X"6D",X"14",X"A1",
		X"49",X"90",X"59",X"61",X"39",X"81",X"38",X"C8",X"20",X"DB",X"6D",X"CF",X"69",X"80",X"31",X"B1",
		X"10",X"BA",X"A1",X"89",X"B0",X"49",X"E3",X"7C",X"32",X"10",X"B6",X"1C",X"65",X"36",X"00",X"07",
		X"C8",X"B8",X"2D",X"CD",X"9E",X"28",X"B5",X"C8",X"D6",X"05",X"B0",X"02",X"B6",X"04",X"6F",X"B6",
		X"23",X"32",X"A2",X"20",X"06",X"8C",X"6D",X"F0",X"95",X"0F",X"8E",X"8B",X"C7",X"22",X"A0",X"20",
		X"45",X"F1",X"CD",X"3C",X"A1",X"B4",X"CD",X"3C",X"A1",X"41",X"26",X"00",X"22",X"00",X"88",X"B4",
		X"65",X"94",X"01",X"B4",X"65",X"94",X"01",X"49",X"18",X"74",X"61",X"B2",X"E8",X"25",X"4F",X"B6",
		X"AC",X"18",X"CB",X"B7",X"4E",X"08",X"26",X"00",X"E7",X"22",X"28",X"88",X"B6",X"10",X"32",X"02",
		X"28",X"45",X"96",X"1E",X"65",X"94",X"01",X"38",X"5B",X"41",X"92",X"69",X"2D",X"6F",X"92",X"68",
		X"8D",X"18",X"6F",X"22",X"28",X"88",X"CD",X"00",X"A1",X"38",X"D3",X"C9",X"4D",X"45",X"A2",X"26",
		X"28",X"6C",X"45",X"A1",X"01",X"F1",X"2C",X"67",X"8A",X"8E",X"28",X"41",X"69",X"C9",X"E3",X"26",
		X"28",X"E7",X"A1",X"B9",X"FE",X"23",X"7E",X"C3",X"C1",X"F4",X"1A",X"48",X"F5",X"1B",X"C9",X"FF",
		X"5F",X"CD",X"75",X"86",X"65",X"65",X"06",X"CD",X"B4",X"87",X"92",X"48",X"B8",X"A7",X"63",X"E7",
		X"48",X"2E",X"29",X"CD",X"89",X"18",X"2E",X"0D",X"39",X"39",X"A6",X"21",X"24",X"8C",X"BA",X"77",
		X"1B",X"23",X"18",X"F2",X"75",X"21",X"80",X"24",X"75",X"36",X"17",X"08",X"89",X"08",X"A0",X"22",
		X"22",X"8C",X"CD",X"1D",X"31",X"2E",X"A8",X"4D",X"AE",X"07",X"4D",X"B6",X"A9",X"18",X"DD",X"77",
		X"A1",X"B6",X"20",X"19",X"75",X"77",X"A0",X"C5",X"43",X"88",X"2C",X"CD",X"6A",X"98",X"88",X"81",
		X"CD",X"8E",X"30",X"20",X"AF",X"CD",X"1F",X"30",X"20",X"0A",X"CD",X"9E",X"30",X"20",X"2D",X"CD",
		X"8D",X"90",X"A0",X"9D",X"65",X"63",X"80",X"2C",X"F1",X"FE",X"A1",X"AF",X"7D",X"D7",X"A2",X"50",
		X"5E",X"89",X"0F",X"75",X"77",X"8B",X"CD",X"CE",X"A6",X"E1",X"AD",X"88",X"95",X"E1",X"38",X"17",
		X"B6",X"4B",X"7D",X"BE",X"17",X"7D",X"D7",X"B7",X"B6",X"98",X"92",X"8A",X"28",X"6D",X"9A",X"A7",
		X"B6",X"A9",X"32",X"8A",X"88",X"65",X"B2",X"A7",X"C9",X"6B",X"6E",X"69",X"28",X"B7",X"F7",X"F7",
		X"57",X"F7",X"57",X"F7",X"57",X"88",X"99",X"CE",X"06",X"FD",X"6D",X"F4",X"05",X"CE",X"A3",X"B1",
		X"7D",X"A6",X"4B",X"2F",X"A5",X"C8",X"30",X"EF",X"30",X"FE",X"30",X"E5",X"30",X"1A",X"B9",X"28",
		X"07",X"00",X"A7",X"16",X"A0",X"92",X"A2",X"28",X"B8",X"8D",X"B6",X"A9",X"92",X"8A",X"28",X"36",
		X"38",X"65",X"09",X"A6",X"BE",X"99",X"CD",X"1A",X"A6",X"61",X"CD",X"09",X"A6",X"65",X"1A",X"A6",
		X"69",X"A1",X"A0",X"89",X"9E",X"BC",X"6D",X"03",X"06",X"A1",X"A0",X"80",X"9E",X"BC",X"6D",X"03",
		X"A6",X"61",X"29",X"88",X"29",X"96",X"20",X"65",X"90",X"A6",X"29",X"BB",X"29",X"96",X"20",X"65",
		X"18",X"A6",X"69",X"FD",X"6D",X"E7",X"01",X"F9",X"D3",X"FD",X"99",X"88",X"A4",X"31",X"B2",X"8A",
		X"88",X"DF",X"59",X"04",X"3D",X"88",X"C4",X"61",X"5D",X"65",X"E7",X"A1",X"59",X"DB",X"5D",X"91",
		X"A0",X"8C",X"B9",X"12",X"A2",X"28",X"D7",X"F9",X"8C",X"B5",X"80",X"64",X"69",X"A6",X"21",X"12",
		X"B9",X"28",X"07",X"08",X"2A",X"86",X"28",X"58",X"32",X"8A",X"88",X"86",X"AF",X"E5",X"AE",X"AD",
		X"4D",X"16",X"27",X"B8",X"0F",X"EE",X"A2",X"E7",X"B6",X"AD",X"19",X"AF",X"4E",X"89",X"EF",X"4D",
		X"6B",X"88",X"88",X"65",X"D6",X"A6",X"49",X"05",X"20",X"46",X"49",X"90",X"40",X"61",X"B6",X"B8",
		X"65",X"94",X"01",X"B4",X"65",X"94",X"01",X"B4",X"65",X"16",X"01",X"CD",X"14",X"81",X"94",X"CD",
		X"B4",X"29",X"B4",X"C9",X"B2",X"19",X"88",X"07",X"C8",X"2E",X"20",X"4D",X"AE",X"00",X"C5",X"6B",
		X"A0",X"20",X"65",X"86",X"07",X"B6",X"A1",X"CD",X"F9",X"80",X"69",X"38",X"4E",X"C9",X"96",X"01",
		X"2E",X"1C",X"4D",X"CD",X"A5",X"29",X"49",X"38",X"D1",X"C9",X"CD",X"84",X"A7",X"CD",X"AA",X"30",
		X"90",X"F0",X"E5",X"6B",X"98",X"25",X"65",X"A1",X"07",X"CD",X"AC",X"87",X"82",X"B8",X"2D",X"78",
		X"F9",X"CD",X"99",X"2D",X"A0",X"F3",X"CD",X"0A",X"30",X"B0",X"C6",X"C5",X"6B",X"B2",X"8D",X"CD",
		X"09",X"87",X"65",X"2C",X"07",X"A2",X"98",X"25",X"58",X"F9",X"65",X"31",X"05",X"A0",X"DB",X"A2",
		X"12",X"8D",X"CD",X"99",X"A5",X"A0",X"C3",X"CD",X"AA",X"30",X"B0",X"E6",X"C5",X"6B",X"14",X"8D",
		X"65",X"A1",X"07",X"C9",X"65",X"3D",X"07",X"0F",X"2F",X"4E",X"A3",X"EF",X"65",X"37",X"07",X"0F",
		X"0F",X"4E",X"2C",X"6F",X"C9",X"CD",X"F4",X"2D",X"46",X"07",X"D6",X"06",X"30",X"F7",X"C9",X"CD",
		X"54",X"85",X"EE",X"0F",X"F6",X"0F",X"98",X"FF",X"61",X"C5",X"4B",X"08",X"28",X"B6",X"34",X"4B",
		X"28",X"2F",X"B2",X"C0",X"8D",X"6F",X"B6",X"0C",X"18",X"CB",X"B7",X"4E",X"A8",X"26",X"28",X"E7",
		X"8A",X"08",X"28",X"B6",X"B6",X"CD",X"14",X"81",X"18",X"F3",X"89",X"69",X"2D",X"2E",X"31",X"87",
		X"77",X"23",X"38",X"FC",X"B2",X"C0",X"8D",X"6F",X"4D",X"CD",X"0C",X"2F",X"60",X"E1",X"39",X"0B",
		X"24",X"CD",X"39",X"85",X"80",X"FB",X"19",X"07",X"24",X"CD",X"39",X"85",X"80",X"E3",X"19",X"03",
		X"38",X"CD",X"99",X"2D",X"A0",X"E3",X"39",X"0F",X"38",X"CD",X"99",X"2D",X"A0",X"DB",X"CD",X"0A",
		X"30",X"B0",X"5E",X"45",X"A5",X"30",X"49",X"38",X"CF",X"41",X"78",X"71",X"B2",X"C0",X"8D",X"6F",
		X"89",X"4A",X"25",X"4D",X"ED",X"EE",X"8B",X"CE",X"C8",X"E1",X"65",X"99",X"0D",X"A0",X"02",X"41",
		X"49",X"AB",X"AB",X"38",X"C6",X"6A",X"63",X"87",X"41",X"C9",X"49",X"BF",X"41",X"B2",X"49",X"8D",
		X"A7",X"9E",X"80",X"FF",X"89",X"4A",X"25",X"B9",X"D9",X"83",X"D8",X"81",X"E1",X"8D",X"9C",X"69",
		X"45",X"8E",X"30",X"40",X"45",X"AC",X"30",X"55",X"BC",X"01",X"45",X"E9",X"30",X"30",X"A5",X"45",
		X"B7",X"30",X"60",X"6D",X"BD",X"30",X"75",X"95",X"81",X"6D",X"FE",X"30",X"10",X"BE",X"65",X"9E",
		X"30",X"40",X"45",X"BC",X"30",X"55",X"BD",X"00",X"45",X"03",X"31",X"30",X"AF",X"45",X"05",X"30",
		X"60",X"6D",X"E3",X"30",X"75",X"94",X"80",X"6D",X"90",X"31",X"10",X"28",X"65",X"8E",X"98",X"48",
		X"45",X"97",X"30",X"48",X"45",X"9E",X"30",X"48",X"45",X"97",X"30",X"48",X"59",X"41",X"C5",X"63",
		X"88",X"8C",X"84",X"6D",X"62",X"30",X"61",X"65",X"43",X"20",X"24",X"8D",X"10",X"55",X"6D",X"EB",
		X"20",X"8C",X"25",X"30",X"C6",X"C5",X"63",X"20",X"8C",X"24",X"30",X"E7",X"C5",X"63",X"20",X"8C",
		X"84",X"6D",X"F2",X"30",X"61",X"65",X"43",X"20",X"24",X"8D",X"10",X"55",X"6D",X"EB",X"88",X"8C",
		X"25",X"30",X"C6",X"C5",X"63",X"20",X"8C",X"24",X"30",X"E7",X"3E",X"46",X"30",X"06",X"3E",X"C6",
		X"10",X"2A",X"96",X"0E",X"89",X"27",X"24",X"F1",X"0F",X"46",X"87",X"8F",X"87",X"8F",X"BA",X"92",
		X"25",X"8C",X"3E",X"00",X"70",X"31",X"4B",X"24",X"8C",X"55",X"BC",X"03",X"45",X"1D",X"31",X"55",
		X"9C",X"2B",X"65",X"BD",X"99",X"69",X"75",X"95",X"83",X"6D",X"15",X"31",X"75",X"95",X"83",X"6D",
		X"35",X"B9",X"61",X"DD",X"9D",X"2A",X"65",X"35",X"B9",X"DD",X"9D",X"2A",X"65",X"35",X"B9",X"C9",
		X"75",X"9C",X"82",X"65",X"15",X"31",X"75",X"9C",X"82",X"65",X"15",X"31",X"61",X"E5",X"43",X"22",
		X"04",X"79",X"2F",X"3C",X"47",X"78",X"2F",X"D6",X"36",X"ED",X"4C",X"47",X"E5",X"43",X"28",X"00",
		X"1E",X"20",X"65",X"B4",X"09",X"65",X"1C",X"A1",X"84",X"E5",X"C3",X"28",X"20",X"65",X"1C",X"A1",
		X"65",X"B4",X"A1",X"DD",X"9C",X"B7",X"92",X"31",X"00",X"A7",X"6C",X"66",X"B9",X"C9",X"96",X"2A",
		X"65",X"59",X"08",X"61",X"7D",X"89",X"88",X"18",X"A7",X"1E",X"80",X"57",X"7D",X"11",X"65",X"F7",
		X"B9",X"28",X"2D",X"7E",X"6E",X"26",X"10",X"2A",X"D6",X"2F",X"F5",X"77",X"28",X"23",X"65",X"F7",
		X"99",X"80",X"85",X"D6",X"E6",X"38",X"10",X"2B",X"5E",X"87",X"1C",X"F5",X"DF",X"29",X"61",X"92",
		X"30",X"00",X"AF",X"C8",X"92",X"3E",X"00",X"E6",X"29",X"C9",X"F5",X"21",X"D8",X"07",X"8B",X"23",
		X"A7",X"1E",X"80",X"57",X"7D",X"11",X"D6",X"92",X"10",X"88",X"AF",X"80",X"91",X"92",X"96",X"88",
		X"EE",X"29",X"80",X"22",X"D2",X"2F",X"EE",X"2B",X"57",X"7A",X"EE",X"D4",X"BB",X"57",X"F5",X"72",
		X"80",X"8B",X"5E",X"F5",X"DF",X"29",X"61",X"89",X"88",X"18",X"86",X"38",X"9E",X"28",X"8B",X"18",
		X"D3",X"C9",X"75",X"21",X"08",X"05",X"75",X"36",X"28",X"F0",X"75",X"36",X"29",X"F8",X"75",X"36",
		X"82",X"A8",X"75",X"9E",X"83",X"AB",X"75",X"9E",X"84",X"29",X"75",X"9E",X"86",X"AA",X"75",X"9E",
		X"2F",X"28",X"75",X"36",X"21",X"28",X"75",X"36",X"36",X"28",X"75",X"36",X"37",X"29",X"61",X"DD",
		X"89",X"28",X"25",X"65",X"04",X"32",X"75",X"89",X"88",X"8D",X"65",X"AC",X"9A",X"75",X"89",X"68",
		X"8D",X"45",X"AC",X"32",X"55",X"A9",X"60",X"8D",X"45",X"0C",X"32",X"41",X"45",X"2F",X"32",X"45",
		X"1A",X"32",X"65",X"EE",X"9A",X"7D",X"5E",X"2E",X"75",X"D7",X"14",X"7D",X"9E",X"2F",X"80",X"7D",
		X"BE",X"08",X"D7",X"55",X"BE",X"09",X"28",X"55",X"BE",X"15",X"D7",X"45",X"E6",X"32",X"41",X"87",
		X"75",X"D7",X"80",X"7D",X"DF",X"29",X"65",X"CE",X"9B",X"69",X"65",X"F4",X"0D",X"46",X"83",X"7D",
		X"FF",X"04",X"45",X"8F",X"A0",X"B5",X"CE",X"07",X"4E",X"01",X"55",X"FF",X"2B",X"41",X"45",X"8F",
		X"08",X"B5",X"63",X"B7",X"63",X"B7",X"C7",X"B2",X"11",X"88",X"AF",X"A0",X"02",X"B2",X"C0",X"18",
		X"A7",X"2F",X"2F",X"CE",X"2B",X"08",X"6F",X"B6",X"AC",X"18",X"55",X"FF",X"2E",X"41",X"55",X"BE",
		X"17",X"AE",X"65",X"8F",X"08",X"76",X"85",X"58",X"75",X"F6",X"85",X"76",X"84",X"48",X"75",X"96",
		X"BF",X"00",X"41",X"55",X"A9",X"A0",X"8D",X"55",X"BE",X"00",X"28",X"55",X"BE",X"01",X"28",X"55",
		X"9E",X"2B",X"01",X"7D",X"9E",X"2E",X"83",X"7D",X"9E",X"2F",X"80",X"7D",X"9E",X"3E",X"80",X"7D",
		X"BE",X"17",X"28",X"55",X"BE",X"1F",X"28",X"45",X"83",X"39",X"41",X"87",X"A9",X"C0",X"8C",X"39",
		X"85",X"28",X"86",X"2D",X"DF",X"B9",X"DF",X"83",X"90",X"D2",X"DF",X"69",X"1A",X"3F",X"20",X"07",
		X"40",X"B2",X"22",X"88",X"CE",X"1F",X"48",X"29",X"29",X"22",X"B2",X"16",X"88",X"43",X"6F",X"A0",
		X"83",X"89",X"93",X"22",X"1A",X"22",X"20",X"6B",X"4F",X"A0",X"07",X"6D",X"74",X"EB",X"9E",X"39",
		X"24",X"45",X"DC",X"4B",X"BE",X"11",X"45",X"F9",X"32",X"41",X"45",X"DC",X"EB",X"BE",X"28",X"24",
		X"65",X"DC",X"43",X"96",X"80",X"6D",X"7D",X"32",X"61",X"B6",X"90",X"B8",X"82",X"B6",X"04",X"86",
		X"28",X"2E",X"20",X"22",X"28",X"00",X"0E",X"24",X"65",X"A5",X"A1",X"10",X"D3",X"C9",X"75",X"21",
		X"80",X"8D",X"10",X"38",X"75",X"89",X"88",X"8D",X"10",X"AA",X"75",X"89",X"C0",X"8D",X"10",X"2C",
		X"75",X"21",X"E8",X"05",X"75",X"7E",X"37",X"11",X"A5",X"BB",X"6B",X"07",X"A5",X"7B",X"BB",X"FF",
		X"9B",X"05",X"9B",X"85",X"1A",X"15",X"19",X"53",X"19",X"E4",X"1A",X"F9",X"9B",X"72",X"9B",X"5F",
		X"B2",X"6E",X"B3",X"F5",X"B3",X"9C",X"B3",X"71",X"BB",X"63",X"B4",X"C3",X"B4",X"E5",X"BB",X"A4",
		X"1D",X"72",X"9B",X"0E",X"85",X"18",X"7E",X"61",X"61",X"75",X"9E",X"28",X"80",X"75",X"9E",X"29",
		X"28",X"CD",X"46",X"BB",X"75",X"34",X"37",X"C9",X"75",X"36",X"37",X"28",X"61",X"DD",X"9E",X"37",
		X"81",X"61",X"75",X"9E",X"17",X"AE",X"61",X"65",X"D7",X"B1",X"75",X"63",X"01",X"6E",X"64",X"0D",
		X"BB",X"CD",X"06",X"BB",X"61",X"DD",X"9E",X"22",X"2C",X"DD",X"9E",X"21",X"27",X"C9",X"92",X"AC",
		X"20",X"AF",X"E0",X"75",X"5E",X"AA",X"1D",X"80",X"84",X"75",X"DF",X"AA",X"61",X"75",X"9E",X"A9",
		X"28",X"DD",X"9C",X"37",X"61",X"CD",X"7F",X"B1",X"75",X"34",X"2F",X"DD",X"D6",X"2F",X"75",X"BE",
		X"86",X"70",X"75",X"9E",X"87",X"28",X"65",X"D8",X"9B",X"89",X"66",X"33",X"ED",X"75",X"5E",X"2C",
		X"19",X"4E",X"BB",X"C3",X"07",X"A5",X"AA",X"B1",X"A4",X"B1",X"BE",X"B1",X"68",X"B1",X"75",X"7E",
		X"85",X"75",X"ED",X"E9",X"65",X"7C",X"99",X"61",X"75",X"D6",X"80",X"EE",X"07",X"F6",X"00",X"68",
		X"75",X"7E",X"29",X"E6",X"27",X"C0",X"92",X"75",X"04",X"FE",X"2A",X"30",X"3E",X"3A",X"10",X"05",
		X"7E",X"2B",X"98",X"B2",X"7E",X"2A",X"88",X"2C",X"2F",X"9A",X"8B",X"88",X"1A",X"23",X"20",X"F6",
		X"2B",X"B0",X"A3",X"55",X"F6",X"1E",X"D6",X"09",X"B8",X"57",X"55",X"BE",X"BC",X"07",X"45",X"7C",
		X"0D",X"46",X"83",X"4E",X"01",X"7D",X"DF",X"BE",X"1E",X"2B",X"9A",X"93",X"24",X"8E",X"7F",X"6D",
		X"89",X"18",X"2E",X"08",X"45",X"89",X"B8",X"2E",X"29",X"45",X"4F",X"18",X"30",X"33",X"45",X"8F",
		X"08",X"B5",X"07",X"AF",X"EE",X"2B",X"E6",X"2B",X"C7",X"B2",X"30",X"8D",X"38",X"90",X"04",X"6D",
		X"EE",X"32",X"5E",X"01",X"55",X"FF",X"BC",X"55",X"BE",X"1E",X"2A",X"B2",X"FD",X"8C",X"D6",X"01",
		X"18",X"AF",X"FD",X"6D",X"46",X"32",X"F6",X"29",X"E1",X"18",X"75",X"D7",X"14",X"7D",X"9E",X"BE",
		X"2A",X"55",X"F6",X"1E",X"39",X"6A",X"34",X"4B",X"8F",X"2D",X"BE",X"35",X"E9",X"36",X"6B",X"38",
		X"22",X"37",X"E2",X"37",X"7A",X"37",X"41",X"36",X"41",X"36",X"7A",X"37",X"24",X"34",X"24",X"34",
		X"8C",X"34",X"8C",X"34",X"58",X"34",X"2B",X"35",X"AC",X"35",X"3D",X"35",X"55",X"F6",X"29",X"D6",
		X"F8",X"A0",X"0C",X"76",X"90",X"A0",X"08",X"7D",X"5E",X"28",X"7E",X"D8",X"08",X"3A",X"7E",X"B8",
		X"A0",X"0E",X"55",X"F6",X"BE",X"5E",X"A9",X"CE",X"2B",X"55",X"FF",X"04",X"45",X"D6",X"B0",X"41",
		X"65",X"F4",X"0D",X"46",X"81",X"7D",X"DF",X"2C",X"E6",X"AD",X"75",X"D7",X"16",X"41",X"61",X"6D",
		X"F4",X"2D",X"CE",X"01",X"4E",X"02",X"55",X"FF",X"2C",X"4E",X"AD",X"55",X"FF",X"1E",X"C9",X"41",
		X"75",X"F6",X"81",X"76",X"90",X"A0",X"14",X"6D",X"58",X"B6",X"75",X"F6",X"84",X"99",X"A9",X"6B",
		X"45",X"8F",X"A5",X"D6",X"BC",X"A0",X"AC",X"D6",X"BD",X"A0",X"A8",X"D6",X"BE",X"A0",X"2C",X"45",
		X"F6",X"B0",X"61",X"7D",X"9E",X"2A",X"60",X"7D",X"9E",X"AB",X"86",X"7D",X"DF",X"BC",X"75",X"96",
		X"37",X"39",X"61",X"DD",X"D6",X"29",X"F6",X"D8",X"80",X"C1",X"10",X"43",X"75",X"7E",X"28",X"FE",
		X"10",X"80",X"E8",X"10",X"E2",X"75",X"5E",X"28",X"7E",X"D8",X"08",X"5F",X"10",X"91",X"65",X"A8",
		X"BE",X"DD",X"46",X"38",X"F5",X"21",X"88",X"05",X"F5",X"7E",X"2C",X"11",X"B9",X"BD",X"6B",X"07",
		X"0D",X"B1",X"9D",X"FD",X"9D",X"73",X"9D",X"89",X"9D",X"0E",X"83",X"63",X"59",X"88",X"06",X"0E",
		X"2A",X"CB",X"D9",X"20",X"20",X"06",X"28",X"CB",X"C9",X"20",X"26",X"06",X"29",X"DD",X"D6",X"35",
		X"75",X"DF",X"16",X"75",X"5E",X"BC",X"75",X"DF",X"86",X"75",X"D8",X"2C",X"61",X"0E",X"82",X"63",
		X"D9",X"20",X"C2",X"06",X"2B",X"CB",X"D1",X"20",X"CC",X"06",X"29",X"CB",X"C1",X"20",X"C2",X"06",
		X"80",X"10",X"72",X"0E",X"80",X"63",X"C9",X"88",X"F4",X"0E",X"81",X"63",X"49",X"88",X"66",X"0E",
		X"2A",X"CB",X"D9",X"20",X"5C",X"06",X"2B",X"18",X"4C",X"06",X"29",X"CB",X"C1",X"20",X"96",X"06",
		X"80",X"63",X"C9",X"88",X"38",X"0E",X"83",X"63",X"59",X"88",X"3E",X"0E",X"82",X"10",X"2E",X"F5",
		X"89",X"88",X"05",X"FD",X"D6",X"2C",X"19",X"84",X"BD",X"C3",X"07",X"A5",X"9C",X"BD",X"50",X"BD",
		X"68",X"35",X"78",X"35",X"7D",X"D6",X"80",X"75",X"3E",X"28",X"E0",X"F5",X"5E",X"29",X"75",X"B6",
		X"29",X"D8",X"75",X"7E",X"36",X"DD",X"DF",X"35",X"75",X"36",X"36",X"28",X"96",X"2D",X"75",X"77",
		X"86",X"75",X"9E",X"2F",X"80",X"E9",X"E9",X"61",X"7D",X"D6",X"80",X"75",X"3E",X"28",X"E0",X"F5",
		X"D6",X"29",X"75",X"BE",X"29",X"D0",X"10",X"52",X"F5",X"7E",X"29",X"DD",X"B6",X"29",X"68",X"FD",
		X"5E",X"28",X"75",X"B6",X"80",X"70",X"10",X"CA",X"7D",X"D6",X"81",X"75",X"3E",X"29",X"E0",X"F5",
		X"F6",X"00",X"55",X"96",X"28",X"58",X"30",X"BA",X"55",X"BE",X"38",X"00",X"45",X"78",X"B6",X"45",
		X"07",X"B1",X"88",X"2F",X"75",X"6B",X"90",X"46",X"75",X"94",X"90",X"6D",X"58",X"B6",X"65",X"3F",
		X"B1",X"A8",X"2F",X"55",X"43",X"10",X"C6",X"55",X"BC",X"10",X"45",X"78",X"B6",X"45",X"BB",X"39",
		X"88",X"2F",X"75",X"6B",X"90",X"56",X"75",X"94",X"90",X"6D",X"58",X"B6",X"65",X"BE",X"19",X"80",
		X"2F",X"55",X"43",X"10",X"D6",X"55",X"BC",X"10",X"41",X"B2",X"97",X"8D",X"D6",X"02",X"44",X"9F",
		X"9D",X"7D",X"5E",X"BC",X"75",X"D7",X"86",X"6D",X"00",X"36",X"75",X"F6",X"90",X"46",X"07",X"99",
		X"65",X"36",X"4B",X"8F",X"A5",X"6F",X"36",X"75",X"36",X"E0",X"36",X"1D",X"37",X"52",X"37",X"55",
		X"9E",X"BE",X"82",X"41",X"61",X"7D",X"5E",X"38",X"86",X"2B",X"87",X"B0",X"82",X"98",X"7B",X"7D",
		X"F8",X"04",X"55",X"BC",X"3D",X"55",X"F6",X"15",X"39",X"8E",X"36",X"4B",X"8F",X"2D",X"1E",X"36",
		X"A8",X"36",X"2A",X"36",X"3E",X"36",X"65",X"F0",X"1E",X"7D",X"D9",X"3E",X"75",X"D0",X"97",X"69",
		X"45",X"78",X"B6",X"55",X"F9",X"18",X"55",X"F8",X"B9",X"41",X"45",X"78",X"B6",X"E1",X"E8",X"55",
		X"56",X"3E",X"75",X"DE",X"97",X"6D",X"31",X"A5",X"60",X"7D",X"9E",X"3D",X"7F",X"69",X"65",X"F0",
		X"B6",X"E1",X"E8",X"55",X"76",X"18",X"55",X"7E",X"B9",X"45",X"99",X"2D",X"A0",X"05",X"55",X"BE",
		X"95",X"D7",X"61",X"7D",X"9E",X"BB",X"82",X"7D",X"9E",X"BE",X"82",X"7D",X"9E",X"3D",X"7F",X"69",
		X"45",X"06",X"37",X"45",X"56",X"36",X"55",X"CD",X"C9",X"39",X"39",X"00",X"31",X"96",X"A8",X"01",
		X"8B",X"F6",X"75",X"D7",X"84",X"69",X"75",X"F6",X"84",X"9E",X"80",X"FF",X"89",X"2A",X"9F",X"B9",
		X"D6",X"C9",X"29",X"28",X"2B",X"2A",X"75",X"7E",X"38",X"06",X"2C",X"0E",X"2B",X"DD",X"ED",X"E1",
		X"91",X"39",X"80",X"11",X"87",X"98",X"82",X"D9",X"8B",X"05",X"90",X"D0",X"61",X"65",X"86",X"37",
		X"65",X"F4",X"A5",X"E6",X"2B",X"FE",X"2B",X"30",X"DF",X"DD",X"ED",X"E1",X"16",X"39",X"2B",X"5F",
		X"96",X"28",X"11",X"D6",X"FD",X"65",X"FE",X"36",X"C7",X"F9",X"38",X"80",X"EB",X"75",X"C6",X"2C",
		X"75",X"77",X"2C",X"B8",X"60",X"DD",X"9E",X"22",X"29",X"DD",X"9E",X"21",X"27",X"DD",X"9E",X"37",
		X"81",X"61",X"65",X"F4",X"0D",X"EE",X"81",X"60",X"7D",X"89",X"A0",X"8D",X"75",X"9E",X"84",X"28",
		X"75",X"7E",X"28",X"FD",X"3E",X"28",X"98",X"2E",X"75",X"CB",X"2C",X"4E",X"E5",X"44",X"4F",X"DD",
		X"5E",X"29",X"7D",X"3E",X"81",X"98",X"86",X"75",X"63",X"2C",X"66",X"E5",X"C4",X"38",X"98",X"2D",
		X"75",X"CB",X"2C",X"46",X"61",X"DD",X"63",X"2C",X"B6",X"C9",X"F5",X"21",X"08",X"05",X"F5",X"7E",
		X"80",X"75",X"3E",X"28",X"08",X"BA",X"65",X"F4",X"0D",X"EE",X"87",X"62",X"41",X"36",X"7D",X"D6",
		X"28",X"D6",X"38",X"DD",X"B6",X"28",X"80",X"20",X"6E",X"A8",X"75",X"BE",X"28",X"C2",X"61",X"BE",
		X"86",X"28",X"7D",X"D6",X"81",X"75",X"3E",X"29",X"18",X"29",X"84",X"75",X"D8",X"2C",X"65",X"5E",
		X"B0",X"C9",X"F5",X"21",X"08",X"05",X"F5",X"7E",X"29",X"DD",X"B6",X"29",X"80",X"32",X"65",X"F4",
		X"0D",X"EE",X"87",X"62",X"41",X"36",X"7D",X"D6",X"81",X"7E",X"90",X"75",X"3E",X"29",X"08",X"A8",
		X"6E",X"A8",X"75",X"BE",X"29",X"C2",X"61",X"BE",X"0E",X"2A",X"F5",X"7E",X"28",X"DD",X"B6",X"28",
		X"18",X"29",X"84",X"75",X"D8",X"2C",X"65",X"5E",X"18",X"61",X"7D",X"89",X"A0",X"8D",X"7D",X"D6",
		X"28",X"55",X"96",X"00",X"A0",X"AA",X"45",X"7C",X"A5",X"CE",X"2F",X"42",X"E9",X"36",X"D5",X"F6",
		X"80",X"5E",X"90",X"7D",X"3E",X"28",X"08",X"98",X"E6",X"20",X"75",X"36",X"80",X"A0",X"B1",X"75",
		X"F6",X"01",X"55",X"96",X"29",X"A0",X"49",X"45",X"F4",X"2D",X"CE",X"07",X"42",X"49",X"36",X"D5",
		X"5E",X"29",X"F6",X"38",X"75",X"36",X"81",X"A0",X"2F",X"4E",X"88",X"7D",X"3E",X"29",X"08",X"80",
		X"4B",X"49",X"36",X"B2",X"97",X"8D",X"D6",X"02",X"44",X"9F",X"35",X"45",X"F4",X"2D",X"CE",X"01",
		X"88",X"62",X"7D",X"81",X"A0",X"8D",X"7D",X"F6",X"81",X"7D",X"3E",X"29",X"88",X"A8",X"65",X"F4",
		X"A5",X"CE",X"2F",X"42",X"E9",X"36",X"D5",X"F6",X"28",X"55",X"96",X"00",X"A0",X"08",X"45",X"7C",
		X"0D",X"46",X"87",X"6A",X"41",X"36",X"7D",X"DE",X"81",X"6D",X"5C",X"A5",X"EE",X"38",X"A2",X"DF",
		X"D5",X"76",X"28",X"45",X"F4",X"2D",X"CE",X"10",X"0B",X"77",X"55",X"BE",X"2C",X"00",X"55",X"F6",
		X"80",X"1B",X"98",X"2E",X"75",X"6B",X"84",X"4E",X"6D",X"CC",X"C7",X"7D",X"5E",X"29",X"B2",X"90",
		X"2E",X"55",X"43",X"04",X"CE",X"C5",X"6C",X"18",X"B8",X"06",X"55",X"43",X"2C",X"CE",X"30",X"04",
		X"75",X"6B",X"84",X"B6",X"75",X"6B",X"13",X"96",X"65",X"5E",X"18",X"7D",X"63",X"BB",X"5E",X"68",
		X"55",X"BD",X"BB",X"55",X"F6",X"1B",X"CE",X"7F",X"48",X"55",X"BE",X"1E",X"29",X"41",X"45",X"7C",
		X"0D",X"46",X"83",X"7D",X"DF",X"2C",X"75",X"F6",X"14",X"7D",X"DF",X"2E",X"65",X"F0",X"1E",X"7D",
		X"F6",X"04",X"39",X"A1",X"6B",X"45",X"8F",X"2D",X"40",X"D6",X"38",X"B0",X"2B",X"D6",X"3E",X"50",
		X"75",X"F6",X"14",X"4E",X"10",X"7D",X"DF",X"2E",X"65",X"F0",X"C3",X"6D",X"4F",X"A1",X"1E",X"BC",
		X"B6",X"28",X"43",X"CD",X"22",X"B8",X"90",X"4E",X"75",X"CB",X"33",X"D6",X"6B",X"4E",X"6A",X"05",
		X"65",X"E7",X"09",X"D6",X"7E",X"20",X"61",X"0C",X"84",X"10",X"FD",X"05",X"10",X"52",X"04",X"04",
		X"10",X"C6",X"75",X"7E",X"29",X"FE",X"39",X"D8",X"75",X"35",X"29",X"C9",X"75",X"7E",X"29",X"FE",
		X"F8",X"78",X"75",X"9C",X"81",X"61",X"75",X"D6",X"80",X"F6",X"11",X"70",X"75",X"9D",X"80",X"61",
		X"75",X"7E",X"28",X"FE",X"50",X"D0",X"75",X"34",X"28",X"C9",X"75",X"7E",X"20",X"A7",X"60",X"3A",
		X"8C",X"88",X"EE",X"BF",X"E0",X"10",X"94",X"75",X"5E",X"A8",X"AF",X"60",X"1A",X"24",X"20",X"EE",
		X"37",X"C0",X"75",X"34",X"24",X"DD",X"D6",X"24",X"EE",X"2B",X"68",X"06",X"28",X"DD",X"D6",X"2D",
		X"7E",X"2D",X"08",X"39",X"86",X"26",X"75",X"D6",X"16",X"F6",X"82",X"80",X"00",X"0E",X"0C",X"F6",
		X"21",X"30",X"2A",X"06",X"3A",X"DD",X"9C",X"24",X"75",X"7E",X"2C",X"FE",X"2B",X"20",X"29",X"3D",
		X"A7",X"75",X"63",X"AC",X"D6",X"88",X"81",X"94",X"A0",X"63",X"8F",X"63",X"8F",X"75",X"DF",X"2A",
		X"75",X"7E",X"2C",X"FE",X"2B",X"20",X"2C",X"DD",X"63",X"2A",X"46",X"DD",X"D6",X"2D",X"75",X"E5",
		X"E9",X"65",X"22",X"31",X"61",X"65",X"F1",X"B1",X"75",X"63",X"01",X"6E",X"64",X"4B",X"19",X"65",
		X"06",X"BB",X"61",X"DD",X"9E",X"22",X"2D",X"DD",X"9E",X"21",X"27",X"06",X"2E",X"CD",X"4F",X"30",
		X"61",X"92",X"8C",X"88",X"EE",X"F7",X"E0",X"96",X"C8",X"75",X"9C",X"AC",X"75",X"63",X"04",X"6E",
		X"88",X"2A",X"96",X"EC",X"75",X"CB",X"2C",X"6E",X"80",X"2A",X"63",X"CF",X"75",X"77",X"2A",X"CD",
		X"2B",X"B1",X"61",X"65",X"F1",X"B1",X"75",X"63",X"01",X"6E",X"64",X"29",X"1A",X"65",X"02",X"B2",
		X"41",X"55",X"BE",X"0A",X"A8",X"55",X"BE",X"09",X"AF",X"41",X"B2",X"24",X"88",X"8F",X"48",X"55",
		X"5E",X"AA",X"1D",X"A0",X"11",X"7D",X"DF",X"AA",X"86",X"A9",X"63",X"CF",X"88",X"A9",X"65",X"8F",
		X"A0",X"B5",X"CE",X"07",X"4E",X"01",X"6F",X"55",X"F8",X"03",X"45",X"AB",X"B1",X"41",X"55",X"F6",
		X"80",X"8E",X"83",X"76",X"10",X"A0",X"13",X"8E",X"82",X"76",X"70",X"A0",X"95",X"7D",X"5E",X"29",
		X"2E",X"01",X"D6",X"10",X"A0",X"0C",X"2E",X"00",X"D6",X"F0",X"A0",X"06",X"45",X"7C",X"A5",X"CE",
		X"83",X"CF",X"75",X"D0",X"84",X"6D",X"27",X"A0",X"1D",X"46",X"87",X"4E",X"81",X"7D",X"DF",X"2B",
		X"45",X"AB",X"B1",X"55",X"BE",X"1E",X"2A",X"55",X"BE",X"1F",X"2A",X"41",X"55",X"43",X"A9",X"46",
		X"64",X"77",X"1A",X"6D",X"B2",X"B2",X"61",X"7D",X"9E",X"AA",X"00",X"7D",X"9E",X"A9",X"07",X"7D",
		X"BE",X"02",X"08",X"45",X"83",X"39",X"39",X"0A",X"28",X"45",X"87",X"28",X"2E",X"02",X"45",X"C7",
		X"10",X"69",X"1A",X"24",X"20",X"07",X"E0",X"7D",X"5E",X"AA",X"1D",X"A0",X"84",X"7D",X"DF",X"AA",
		X"41",X"55",X"BE",X"09",X"28",X"55",X"BC",X"1F",X"A9",X"98",X"8D",X"BD",X"41",X"55",X"BC",X"07",
		X"75",X"F6",X"87",X"7D",X"3E",X"2E",X"70",X"7D",X"9E",X"2F",X"80",X"7D",X"5E",X"28",X"EE",X"AF",
		X"D6",X"08",X"A8",X"0F",X"55",X"F6",X"29",X"CE",X"AF",X"A8",X"A8",X"55",X"BE",X"09",X"28",X"55",
		X"9C",X"BF",X"61",X"6D",X"39",X"33",X"61",X"65",X"43",X"00",X"25",X"B2",X"AC",X"8D",X"91",X"A2",
		X"B3",X"45",X"8F",X"2D",X"55",X"F9",X"28",X"55",X"F8",X"01",X"B2",X"A4",X"8D",X"55",X"FF",X"04",
		X"EE",X"2A",X"C7",X"B2",X"AC",X"8D",X"0F",X"46",X"81",X"10",X"7E",X"2B",X"88",X"29",X"1D",X"0F",
		X"6E",X"3A",X"0F",X"07",X"75",X"77",X"2A",X"DD",X"D6",X"2C",X"F6",X"2A",X"88",X"2C",X"75",X"CB",
		X"82",X"CE",X"75",X"9E",X"86",X"2B",X"1A",X"07",X"25",X"75",X"DF",X"2F",X"65",X"CE",X"9B",X"65",
		X"83",X"B1",X"75",X"36",X"21",X"28",X"75",X"34",X"37",X"C9",X"BA",X"B3",X"BF",X"B3",X"B4",X"B3",
		X"C1",X"B3",X"58",X"7E",X"90",X"4F",X"61",X"D0",X"E6",X"38",X"C7",X"61",X"59",X"7E",X"90",X"47",
		X"61",X"79",X"6E",X"38",X"47",X"C9",X"75",X"7E",X"20",X"A7",X"80",X"3A",X"75",X"34",X"2F",X"DD",
		X"5E",X"2F",X"75",X"B6",X"86",X"70",X"75",X"9E",X"87",X"28",X"65",X"91",X"9B",X"61",X"75",X"D6",
		X"2C",X"FE",X"2B",X"20",X"29",X"3D",X"2F",X"C6",X"24",X"07",X"0F",X"DD",X"DF",X"2A",X"75",X"7E",
		X"84",X"F6",X"83",X"88",X"84",X"75",X"63",X"2A",X"66",X"65",X"2B",X"B1",X"61",X"75",X"63",X"A9",
		X"6E",X"CC",X"00",X"B3",X"65",X"06",X"BB",X"C9",X"75",X"36",X"22",X"29",X"75",X"36",X"21",X"27",
		X"75",X"D6",X"84",X"F6",X"83",X"88",X"81",X"95",X"A7",X"94",X"E6",X"AC",X"87",X"0F",X"75",X"DF",
		X"2A",X"DD",X"D6",X"2C",X"F6",X"2B",X"88",X"2C",X"75",X"CB",X"2A",X"46",X"65",X"83",X"B1",X"DD",
		X"9E",X"A8",X"7F",X"61",X"75",X"63",X"01",X"6E",X"64",X"97",X"1B",X"65",X"8A",X"B4",X"61",X"75",
		X"9E",X"22",X"2C",X"DD",X"9E",X"21",X"27",X"DD",X"D6",X"32",X"AF",X"20",X"24",X"DD",X"9E",X"28",
		X"80",X"75",X"9E",X"29",X"80",X"65",X"66",X"33",X"61",X"65",X"6E",X"B3",X"65",X"A9",X"1C",X"75",
		X"9C",X"28",X"75",X"34",X"29",X"CD",X"F0",X"B6",X"96",X"3B",X"65",X"4C",X"63",X"C9",X"75",X"7E",
		X"12",X"95",X"A7",X"1E",X"80",X"57",X"89",X"29",X"1C",X"11",X"56",X"8B",X"D6",X"65",X"2F",X"A0",
		X"41",X"28",X"28",X"A0",X"28",X"40",X"29",X"80",X"2A",X"55",X"F6",X"1A",X"CE",X"07",X"B5",X"3E",
		X"80",X"FF",X"89",X"BE",X"1C",X"B9",X"5E",X"7D",X"DF",X"2A",X"65",X"83",X"19",X"69",X"A4",X"88",
		X"8C",X"90",X"B2",X"24",X"88",X"8F",X"48",X"55",X"F6",X"0A",X"B5",X"A0",X"2C",X"55",X"FF",X"0A",
		X"61",X"7D",X"9E",X"A9",X"80",X"7D",X"9C",X"BF",X"65",X"F0",X"1E",X"6D",X"70",X"EB",X"89",X"98",
		X"8D",X"BD",X"A9",X"DF",X"8D",X"BE",X"08",X"A3",X"BE",X"08",X"41",X"A9",X"DD",X"8D",X"F6",X"8F",
		X"88",X"BA",X"75",X"96",X"17",X"28",X"65",X"8F",X"08",X"B5",X"07",X"AF",X"EE",X"2B",X"E6",X"2C",
		X"6F",X"B2",X"98",X"8D",X"90",X"58",X"B6",X"04",X"BA",X"BB",X"8C",X"41",X"BD",X"A9",X"4A",X"8D",
		X"46",X"83",X"C6",X"83",X"58",X"09",X"08",X"D0",X"E5",X"6D",X"E6",X"6A",X"E1",X"6D",X"76",X"B4",
		X"55",X"F9",X"28",X"55",X"F8",X"01",X"45",X"CE",X"33",X"55",X"BE",X"02",X"DC",X"45",X"8F",X"28",
		X"1D",X"46",X"87",X"B4",X"75",X"D7",X"83",X"6D",X"2B",X"B1",X"75",X"F6",X"14",X"7D",X"DF",X"2E",
		X"55",X"BE",X"A9",X"00",X"55",X"BE",X"AB",X"06",X"45",X"7C",X"A5",X"CE",X"2F",X"B4",X"55",X"FF",
		X"16",X"7D",X"9E",X"BB",X"94",X"7D",X"9C",X"BF",X"86",X"2B",X"65",X"4F",X"10",X"81",X"16",X"8D",
		X"39",X"20",X"28",X"2E",X"2C",X"B6",X"2A",X"96",X"40",X"31",X"38",X"FB",X"A9",X"1F",X"8D",X"2E",
		X"84",X"B6",X"82",X"36",X"08",X"2C",X"11",X"98",X"7A",X"69",X"0B",X"96",X"82",X"69",X"58",X"8F",
		X"2F",X"2F",X"6F",X"F1",X"4E",X"02",X"2F",X"2F",X"2F",X"67",X"41",X"55",X"43",X"09",X"6E",X"44",
		X"FE",X"B4",X"65",X"D7",X"1C",X"69",X"75",X"96",X"02",X"2C",X"75",X"96",X"01",X"AF",X"61",X"B2",
		X"AC",X"00",X"EE",X"B7",X"68",X"DD",X"D6",X"22",X"95",X"28",X"2C",X"DD",X"DF",X"22",X"61",X"DD",
		X"5E",X"AB",X"1D",X"80",X"93",X"75",X"DF",X"AB",X"75",X"9E",X"01",X"28",X"75",X"D6",X"82",X"7E",
		X"2C",X"DD",X"DF",X"2A",X"65",X"83",X"B1",X"C9",X"75",X"34",X"37",X"C9",X"75",X"CB",X"21",X"6E",
		X"64",X"56",X"1C",X"65",X"9F",X"B5",X"61",X"92",X"8C",X"88",X"EE",X"B7",X"E0",X"75",X"5E",X"AA",
		X"95",X"28",X"2C",X"DD",X"DF",X"22",X"61",X"DD",X"D6",X"23",X"95",X"28",X"3B",X"DD",X"DF",X"23",
		X"75",X"9E",X"01",X"28",X"75",X"D6",X"82",X"6E",X"84",X"75",X"DF",X"2A",X"65",X"83",X"19",X"61",
		X"75",X"34",X"37",X"21",X"10",X"05",X"9D",X"DD",X"9E",X"28",X"28",X"DD",X"9E",X"29",X"28",X"CD",
		X"66",X"33",X"61",X"75",X"89",X"08",X"25",X"75",X"5E",X"BF",X"91",X"08",X"1D",X"6B",X"27",X"A5",
		X"70",X"BB",X"18",X"B5",X"97",X"B5",X"C1",X"B7",X"7B",X"68",X"12",X"68",X"9B",X"B7",X"E0",X"BB",
		X"65",X"EA",X"19",X"75",X"63",X"A9",X"C6",X"64",X"36",X"B5",X"65",X"07",X"1D",X"61",X"75",X"9E",
		X"22",X"2A",X"75",X"36",X"21",X"27",X"61",X"3A",X"AC",X"00",X"AF",X"C0",X"75",X"7E",X"22",X"3D",
		X"08",X"2C",X"75",X"DF",X"02",X"61",X"75",X"9E",X"01",X"28",X"75",X"9E",X"17",X"2A",X"61",X"75",
		X"89",X"08",X"05",X"CD",X"62",X"B1",X"75",X"34",X"2F",X"DD",X"D6",X"2F",X"75",X"BE",X"2E",X"D8",
		X"75",X"9E",X"87",X"28",X"65",X"2E",X"1E",X"89",X"EC",X"B5",X"ED",X"75",X"5E",X"2C",X"91",X"C6",
		X"B5",X"C3",X"07",X"A5",X"75",X"7E",X"2D",X"DD",X"ED",X"E1",X"65",X"7C",X"B9",X"C9",X"DE",X"B5",
		X"7A",X"B5",X"7E",X"B5",X"82",X"B6",X"75",X"9D",X"81",X"61",X"75",X"9C",X"81",X"61",X"75",X"9D",
		X"28",X"41",X"55",X"BC",X"28",X"41",X"55",X"F6",X"28",X"CE",X"AF",X"D6",X"A8",X"A8",X"2F",X"55",
		X"5E",X"29",X"EE",X"AF",X"08",X"2C",X"65",X"06",X"1E",X"69",X"65",X"54",X"1E",X"6D",X"A0",X"B7",
		X"55",X"43",X"A8",X"46",X"42",X"5C",X"B6",X"45",X"F0",X"3E",X"55",X"F6",X"2C",X"39",X"36",X"3E",
		X"65",X"8F",X"0D",X"68",X"E9",X"69",X"1E",X"B6",X"56",X"B6",X"CF",X"B6",X"4F",X"B6",X"85",X"6D",
		X"6C",X"3E",X"48",X"24",X"45",X"6F",X"A1",X"F6",X"D6",X"20",X"40",X"D6",X"08",X"50",X"D6",X"90",
		X"18",X"A8",X"7E",X"98",X"70",X"76",X"34",X"B0",X"81",X"69",X"3F",X"69",X"E9",X"69",X"84",X"8C",
		X"45",X"44",X"B6",X"48",X"24",X"30",X"DD",X"25",X"45",X"44",X"B6",X"48",X"2C",X"30",X"5D",X"24",
		X"04",X"6D",X"C4",X"B6",X"E0",X"8C",X"10",X"CC",X"75",X"F6",X"80",X"6B",X"1F",X"6B",X"1F",X"6B",
		X"B7",X"5E",X"2A",X"67",X"55",X"F6",X"29",X"43",X"B7",X"43",X"B7",X"43",X"B7",X"6F",X"41",X"D5",
		X"5E",X"28",X"63",X"B7",X"63",X"B7",X"63",X"B7",X"F6",X"2A",X"47",X"75",X"5E",X"29",X"63",X"B7",
		X"43",X"B7",X"43",X"B7",X"6F",X"41",X"B2",X"19",X"88",X"8F",X"40",X"45",X"D3",X"2A",X"A7",X"CE",
		X"07",X"68",X"86",X"2C",X"07",X"B0",X"83",X"98",X"7B",X"69",X"1E",X"2C",X"B0",X"7D",X"3E",X"2C",
		X"40",X"55",X"F6",X"00",X"CE",X"0F",X"D6",X"08",X"A0",X"12",X"D6",X"04",X"50",X"D6",X"AC",X"58",
		X"86",X"2B",X"7E",X"A8",X"18",X"2A",X"86",X"2A",X"75",X"D0",X"84",X"69",X"75",X"F6",X"81",X"46",
		X"AF",X"D6",X"2C",X"B0",X"2B",X"D6",X"AC",X"50",X"2E",X"01",X"D6",X"08",X"B8",X"02",X"2E",X"00",
		X"75",X"D0",X"84",X"69",X"1A",X"B9",X"20",X"07",X"08",X"A5",X"2F",X"92",X"FC",X"8C",X"75",X"96",
		X"20",X"28",X"65",X"D3",X"A2",X"2F",X"EE",X"27",X"60",X"DD",X"9E",X"20",X"D7",X"DD",X"4E",X"2C",
		X"75",X"D8",X"90",X"0E",X"84",X"07",X"18",X"2B",X"90",X"D3",X"61",X"96",X"84",X"38",X"75",X"DF",
		X"2C",X"CB",X"77",X"32",X"DC",X"04",X"61",X"2A",X"DA",X"04",X"19",X"DD",X"04",X"EB",X"12",X"CB",
		X"C6",X"80",X"01",X"1B",X"6D",X"5B",X"FA",X"8C",X"07",X"07",X"07",X"07",X"9C",X"E3",X"63",X"5F",
		X"FD",X"C4",X"13",X"B7",X"F9",X"DD",X"9E",X"20",X"28",X"CB",X"57",X"C8",X"EE",X"2B",X"75",X"77",
		X"84",X"75",X"9E",X"A8",X"7F",X"61",X"65",X"D2",X"1E",X"65",X"A5",X"B7",X"0A",X"52",X"24",X"19",
		X"DD",X"04",X"E3",X"3A",X"DC",X"04",X"63",X"46",X"80",X"3B",X"07",X"0F",X"07",X"0F",X"EE",X"D8",
		X"C7",X"12",X"EE",X"AF",X"B8",X"1A",X"93",X"E5",X"D3",X"52",X"24",X"9C",X"61",X"1A",X"9C",X"61",
		X"92",X"31",X"00",X"A7",X"60",X"CD",X"D3",X"A2",X"87",X"CB",X"D7",X"28",X"A9",X"DD",X"D6",X"27",
		X"1C",X"60",X"75",X"9E",X"07",X"D7",X"89",X"54",X"24",X"63",X"F6",X"92",X"3F",X"8D",X"AF",X"68",
		X"96",X"29",X"9A",X"97",X"05",X"DD",X"9E",X"37",X"2B",X"DD",X"9E",X"23",X"28",X"C9",X"75",X"36",
		X"07",X"28",X"61",X"96",X"16",X"65",X"F1",X"A0",X"65",X"DA",X"1F",X"0E",X"04",X"06",X"12",X"6D",
		X"63",X"40",X"80",X"29",X"04",X"79",X"0F",X"07",X"75",X"77",X"2A",X"CD",X"83",X"B1",X"96",X"20",
		X"65",X"59",X"08",X"69",X"90",X"C1",X"75",X"9C",X"17",X"61",X"2F",X"89",X"FB",X"8F",X"91",X"2A",
		X"28",X"77",X"11",X"77",X"11",X"77",X"11",X"77",X"61",X"DD",X"D6",X"23",X"19",X"DA",X"B7",X"C3",
		X"27",X"A5",X"7A",X"B7",X"8B",X"68",X"17",X"68",X"46",X"68",X"86",X"28",X"75",X"D6",X"84",X"F6");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
