library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"F7",X"F0",X"11",X"11",X"11",X"33",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"F0",X"F7",X"CF",X"C7",X"F0",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"D5",X"91",X"11",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"C0",X"88",X"88",X"88",X"00",
		X"88",X"CC",X"66",X"B3",X"B3",X"C4",X"80",X"B3",X"11",X"CC",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",
		X"F7",X"E6",X"F0",X"E6",X"F7",X"F0",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",
		X"0F",X"09",X"06",X"06",X"06",X"0F",X"00",X"F0",X"07",X"05",X"05",X"05",X"04",X"07",X"00",X"00",
		X"91",X"F7",X"80",X"F7",X"91",X"11",X"88",X"00",X"F0",X"F0",X"FC",X"F0",X"F0",X"F0",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"91",X"08",X"08",X"08",X"08",X"08",X"4F",X"CC",X"F0",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"03",X"03",X"0F",X"0F",X"0F",X"0F",X"03",X"03",
		X"0C",X"0C",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"03",X"03",X"0F",X"0F",X"0F",X"0F",X"00",X"00",
		X"D1",X"D1",X"F3",X"C0",X"F3",X"D1",X"D1",X"CC",X"70",X"F6",X"D4",X"F1",X"D4",X"F6",X"70",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"88",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"00",
		X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"75",X"FA",X"75",X"FA",X"75",X"FA",X"75",X"FA",
		X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"AA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",X"AA",
		X"00",X"EA",X"F5",X"FA",X"F5",X"FA",X"F5",X"EA",X"F5",X"FA",X"F5",X"FA",X"F5",X"FA",X"75",X"00",
		X"EA",X"F5",X"FA",X"F5",X"FA",X"F5",X"EA",X"00",X"00",X"75",X"FA",X"F5",X"FA",X"F5",X"FA",X"F5",
		X"C4",X"EA",X"E4",X"EA",X"F5",X"FA",X"F5",X"EA",X"75",X"FA",X"F5",X"FA",X"75",X"72",X"75",X"32",
		X"EA",X"F5",X"FA",X"F5",X"EA",X"E4",X"EA",X"C4",X"32",X"75",X"72",X"75",X"FA",X"F5",X"FA",X"75",
		X"0C",X"86",X"C3",X"E1",X"E1",X"E9",X"E8",X"C0",X"03",X"70",X"F0",X"F0",X"F4",X"F5",X"71",X"30",
		X"00",X"22",X"44",X"00",X"33",X"00",X"44",X"22",X"00",X"22",X"11",X"00",X"66",X"00",X"11",X"22",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F6",X"F3",X"70",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"21",X"70",X"F3",X"F4",X"F4",X"F0",X"F0",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"E5",X"F4",X"E8",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F0",
		X"0E",X"C3",X"E9",X"ED",X"E5",X"E5",X"E1",X"E1",X"0F",X"F0",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"F8",X"FC",X"FE",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"77",
		X"0F",X"FE",X"FC",X"F8",X"F0",X"0F",X"0F",X"0F",X"03",X"77",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"E1",X"E3",X"E7",X"EF",X"EF",X"EF",X"EE",X"CC",X"1E",X"1E",X"1E",X"1E",X"F1",X"F3",X"F7",X"FF",
		X"0E",X"CF",X"EF",X"EF",X"EF",X"EF",X"E7",X"E3",X"0F",X"FF",X"F7",X"F3",X"F1",X"1E",X"1E",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"EE",X"CC",X"EE",X"FF",X"00",X"00",X"33",X"33",X"77",X"FF",X"77",X"33",X"33",
		X"00",X"0E",X"01",X"0A",X"0C",X"08",X"08",X"0E",X"00",X"03",X"04",X"09",X"0A",X"0A",X"0A",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",
		X"89",X"98",X"F6",X"F0",X"01",X"01",X"01",X"03",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"F0",X"F6",X"98",X"81",X"E1",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"8D",X"81",X"01",X"00",X"00",X"00",X"00",X"00",X"7F",X"7B",X"F0",X"C0",X"08",X"08",X"08",X"00",
		X"08",X"0C",X"06",X"83",X"8B",X"8C",X"88",X"8B",X"01",X"0C",X"F0",X"F3",X"F7",X"7F",X"7F",X"7F",
		X"98",X"F6",X"F0",X"01",X"01",X"01",X"03",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"F0",X"F6",X"98",X"89",X"E1",X"89",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"30",
		X"8D",X"81",X"01",X"00",X"00",X"00",X"00",X"00",X"7F",X"F3",X"F0",X"08",X"08",X"08",X"00",X"00",
		X"01",X"01",X"01",X"83",X"8B",X"8C",X"88",X"8B",X"00",X"0C",X"F0",X"F3",X"7F",X"7F",X"7F",X"7F",
		X"C4",X"C4",X"F2",X"F0",X"70",X"10",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"10",X"34",X"79",X"78",X"E1",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"84",X"86",X"84",X"0C",X"08",X"00",X"00",X"1E",X"90",X"91",X"FE",X"F0",X"E0",X"07",X"00",
		X"0C",X"06",X"06",X"8C",X"CC",X"EC",X"EC",X"E8",X"0E",X"04",X"F7",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"00",X"EE",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"11",X"00",X"00",X"00",
		X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"00",
		X"CC",X"22",X"55",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"AA",X"AA",X"AA",X"99",X"44",X"33",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"0E",X"0C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",X"0E",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0C",X"0E",X"02",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"0E",X"01",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"09",X"0F",X"0F",X"0F",X"07",
		X"00",X"0F",X"0F",X"0F",X"0F",X"02",X"0D",X"0E",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"06",X"0A",X"0E",X"0E",X"0E",X"0E",X"0C",X"01",X"0F",X"0F",X"0F",X"07",X"07",X"0B",X"0F",
		X"00",X"0C",X"0E",X"0E",X"0E",X"0A",X"06",X"0E",X"00",X"0F",X"0B",X"0B",X"07",X"0F",X"0F",X"0E",
		X"0E",X"01",X"0E",X"0E",X"0F",X"07",X"0F",X"0F",X"0E",X"0F",X"0E",X"09",X"0E",X"0F",X"0D",X"07",
		X"00",X"0F",X"0D",X"0F",X"0F",X"02",X"0D",X"0E",X"00",X"07",X"0B",X"0E",X"0F",X"0F",X"0F",X"09",
		X"0E",X"06",X"0A",X"0E",X"0E",X"0E",X"06",X"0C",X"01",X"0F",X"0E",X"0F",X"05",X"07",X"0B",X"0F",
		X"00",X"0C",X"0A",X"0E",X"0E",X"0A",X"06",X"0E",X"00",X"0F",X"0B",X"0B",X"05",X"0F",X"0F",X"0E",
		X"0E",X"01",X"0E",X"0E",X"0D",X"03",X"0F",X"0F",X"06",X"0F",X"0E",X"09",X"06",X"0E",X"0D",X"05",
		X"00",X"0E",X"01",X"0F",X"07",X"02",X"0D",X"0E",X"00",X"07",X"0B",X"08",X"0F",X"0F",X"0E",X"09",
		X"0E",X"06",X"08",X"0E",X"0E",X"0E",X"02",X"0C",X"00",X"0F",X"0E",X"0E",X"05",X"04",X"0B",X"07",
		X"00",X"0C",X"0A",X"0A",X"06",X"0A",X"04",X"0E",X"00",X"0D",X"0B",X"09",X"04",X"0F",X"0F",X"0E",
		X"06",X"00",X"06",X"07",X"06",X"00",X"0D",X"05",X"06",X"0D",X"09",X"00",X"03",X"04",X"06",X"02",
		X"0A",X"0C",X"01",X"07",X"05",X"01",X"06",X"0F",X"00",X"03",X"01",X"04",X"0B",X"0D",X"0E",X"00",
		X"05",X"0B",X"00",X"07",X"06",X"01",X"09",X"0C",X"00",X"03",X"0D",X"06",X"02",X"08",X"09",X"03",
		X"00",X"06",X"08",X"09",X"03",X"0D",X"08",X"06",X"02",X"04",X"01",X"08",X"02",X"06",X"05",X"04",
		X"01",X"04",X"0F",X"01",X"0B",X"00",X"0A",X"0E",X"01",X"03",X"02",X"00",X"01",X"00",X"01",X"00",
		X"02",X"0D",X"04",X"01",X"0D",X"04",X"09",X"03",X"00",X"00",X"00",X"01",X"02",X"01",X"03",X"00",
		X"03",X"0D",X"08",X"07",X"0B",X"01",X"0C",X"0B",X"08",X"01",X"06",X"0A",X"01",X"04",X"0C",X"09",
		X"08",X"01",X"04",X"05",X"0B",X"0B",X"04",X"03",X"08",X"01",X"04",X"0A",X"04",X"04",X"09",X"05",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"0A",X"01",X"03",X"00",X"0D",X"0A",X"0B",X"08",X"02",X"01",X"05",X"00",X"0A",X"04",
		X"02",X"08",X"02",X"0B",X"01",X"05",X"02",X"08",X"00",X"02",X"0A",X"01",X"05",X"08",X"0A",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"02",X"00",X"05",X"01",X"08",X"02",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",
		X"08",X"01",X"00",X"0A",X"00",X"05",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"01",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"02",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F8",X"FB",X"F3",X"F0",X"30",X"00",X"70",X"71",X"31",X"30",X"10",X"00",X"00",X"00",
		X"00",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FC",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"D2",X"2D",X"F8",X"3D",X"D7",X"F0",X"30",X"00",X"25",X"71",X"21",X"30",X"10",X"00",X"00",X"00",
		X"00",X"30",X"F0",X"F0",X"B4",X"78",X"87",X"78",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"52",
		X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"F0",X"F0",X"3C",X"FC",X"F8",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"00",X"C0",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",
		X"D2",X"2D",X"F8",X"3D",X"D7",X"E1",X"21",X"00",X"25",X"71",X"21",X"30",X"01",X"00",X"00",X"00",
		X"00",X"30",X"D2",X"A5",X"78",X"78",X"87",X"78",X"00",X"00",X"00",X"01",X"30",X"30",X"70",X"52",
		X"E0",X"68",X"C0",X"C0",X"80",X"00",X"00",X"00",X"E1",X"D2",X"3C",X"DE",X"69",X"F0",X"C0",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"C2",X"2C",X"00",X"C0",X"D2",X"B4",X"5A",X"69",X"F0",X"3C",
		X"00",X"20",X"D0",X"34",X"DE",X"E5",X"D0",X"30",X"00",X"00",X"00",X"30",X"10",X"10",X"00",X"00",
		X"30",X"F0",X"52",X"B4",X"B0",X"40",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"00",X"00",X"00",
		X"E0",X"60",X"E0",X"68",X"80",X"C0",X"80",X"00",X"20",X"50",X"30",X"D2",X"69",X"BE",X"DC",X"E0",
		X"00",X"80",X"80",X"48",X"E0",X"60",X"E0",X"20",X"60",X"B4",X"5A",X"B4",X"43",X"70",X"A0",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"C3",X"C3",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"C0",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"33",X"FF",X"33",X"33",X"33",X"33",X"33",X"11",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"77",X"00",X"99",X"AA",X"AA",X"AA",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"88",X"77",X"00",X"77",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"11",X"11",X"11",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"11",X"11",X"EE",X"00",X"EE",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"0E",X"0C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"06",X"06",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"01",X"01",X"01",X"12",X"12",X"12",X"12",X"01",
		X"F0",X"F0",X"78",X"78",X"78",X"78",X"78",X"F0",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"34",X"34",X"34",X"34",X"12",X"12",X"12",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"01",X"12",X"34",X"34",X"34",X"78",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"E1",X"86",X"08",X"00",X"00",X"00",X"00",X"F1",X"F0",X"F0",X"E1",X"C2",X"84",X"08",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F3",X"F7",X"FF",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"96",X"09",X"00",X"00",X"00",X"08",X"09",X"96",X"F0",X"F0",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"01",X"1E",X"F0",X"F0",
		X"34",X"34",X"34",X"34",X"12",X"12",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"12",X"12",X"12",X"12",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"FF",X"F8",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"F3",X"7B",X"78",X"78",X"78",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"FE",
		X"34",X"34",X"12",X"12",X"12",X"1A",X"96",X"E1",X"00",X"00",X"00",X"00",X"08",X"87",X"F0",X"F0",
		X"01",X"12",X"12",X"12",X"12",X"34",X"34",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"35",X"35",X"34",X"12",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"16",X"69",X"78",X"78",X"78",X"79",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FE",X"FE",X"F6",X"F7",X"F3",X"78",X"35",X"35",X"34",X"12",X"12",X"01",X"01",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"12",X"12",X"34",X"34",X"34",X"34",X"35",X"35",
		X"F6",X"F7",X"F3",X"79",X"34",X"16",X"69",X"F0",X"12",X"12",X"01",X"00",X"00",X"00",X"00",X"01",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FC",X"78",X"78",X"78",X"78",X"78",X"34",X"34",X"34",
		X"F0",X"78",X"1E",X"E1",X"F0",X"F0",X"F0",X"F0",X"C3",X"E1",X"F0",X"F8",X"FC",X"FE",X"F6",X"7A",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"34",X"34",X"1E",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"F7",X"F6",X"F6",X"F6",X"F2",X"F0",X"F0",
		X"00",X"03",X"3C",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"00",X"00",X"01",X"12",X"34",X"79",X"7B",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"E1",X"D2",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"78",X"B4",X"B4",X"D2",X"D2",X"78",X"96",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"F3",X"F6",X"F6",X"F4",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"87",X"78",X"F0",X"F0",X"FC",X"FE",X"FF",X"FF",X"F0",X"E1",X"1E",X"78",X"F1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",
		X"F0",X"F0",X"F0",X"FC",X"FC",X"F0",X"F0",X"0F",X"F0",X"F0",X"FF",X"FF",X"F7",X"F0",X"78",X"87",
		X"F0",X"F0",X"78",X"78",X"78",X"F0",X"F0",X"F0",X"96",X"09",X"08",X"08",X"84",X"C3",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"96",X"E1",X"F0",X"F0",
		X"34",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"84",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F6",X"F7",X"7B",X"34",X"F0",X"F0",X"F0",X"F0",X"F0",X"C3",X"84",X"08",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"07",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"3C",X"03",X"00",X"00",X"00",X"F0",X"F0",X"1E",X"01",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F3",X"F0",X"3C",X"03",X"00",X"0F",X"F0",X"78",X"16",X"01",X"00",X"00",X"00",X"0F",
		X"FC",X"FE",X"F6",X"F6",X"78",X"78",X"78",X"F0",X"F0",X"96",X"09",X"09",X"08",X"08",X"84",X"C3",
		X"F0",X"F0",X"F0",X"E1",X"1E",X"C3",X"E1",X"F0",X"F0",X"F0",X"F0",X"1E",X"E1",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F7",X"FF",X"F8",X"E1",X"D2",
		X"F0",X"78",X"7B",X"7B",X"7B",X"B5",X"D2",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"D2",X"3C",
		X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"FF",X"FF",X"FE",X"F0",X"E1",X"1E",X"D2",X"F0",X"F0",X"F7",X"F3",X"F0",X"F0",X"0F",X"F0",
		X"08",X"87",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"FF",X"FF",X"FF",X"F0",X"F0",X"0F",X"00",X"FF",X"F7",X"F3",X"F0",X"78",X"07",X"00",X"00",
		X"F1",X"FF",X"FF",X"FF",X"F0",X"C3",X"0C",X"0F",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"0F",X"0F",
		X"D2",X"D2",X"D2",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"B4",X"B4",X"B4",X"D2",X"D2",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F1",X"78",X"96",X"E1",X"F0",X"F0",X"F0",X"F0",X"1E",X"E1",X"F0",X"F0",X"78",
		X"F0",X"F0",X"F0",X"F0",X"F1",X"F0",X"78",X"87",X"F0",X"F0",X"F0",X"F0",X"FE",X"F0",X"0F",X"F0",
		X"B4",X"D2",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"B4",X"B4",X"79",X"79",X"78",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"F0",X"0F",
		X"E1",X"D2",X"B4",X"78",X"F0",X"F0",X"F0",X"F0",X"FF",X"FE",X"F8",X"F0",X"C3",X"3C",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F3",X"F7",
		X"00",X"00",X"00",X"08",X"84",X"C2",X"E1",X"E1",X"00",X"08",X"86",X"E1",X"F0",X"F0",X"F0",X"F0",
		X"F7",X"FF",X"FF",X"FF",X"FC",X"F0",X"F0",X"0F",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"0F",
		X"0E",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E9",X"C2",X"84",X"08",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FC",X"F0",X"87",X"08",X"00",X"0F",
		X"00",X"00",X"08",X"84",X"C2",X"E1",X"E1",X"E1",X"C2",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"ED",X"ED",X"E9",X"E1",X"C2",X"0C",X"00",X"00",X"F0",X"F1",X"FF",X"FF",X"F0",X"C3",X"0C",X"84",
		X"08",X"84",X"C2",X"C2",X"C2",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"CA",X"CA",X"CA",X"CA",X"C2",X"84",X"08",X"00",X"F1",X"F3",X"F7",X"FF",X"FE",X"F0",X"E1",X"0F",
		X"FF",X"FE",X"F0",X"0F",X"84",X"84",X"C2",X"C2",X"F7",X"F1",X"78",X"87",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"84",X"08",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"84",X"84",X"84",X"84",
		X"C2",X"C2",X"84",X"08",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"E1",X"C2",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"08",X"84",X"C2",X"C2",X"00",X"08",X"86",X"E1",X"F0",X"F0",X"F0",X"F0",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"E1",X"86",X"08",X"00",X"00",X"00",X"00",
		X"E1",X"E1",X"E1",X"E1",X"C2",X"C2",X"C2",X"84",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"08",X"84",X"C2",X"E1",X"E1",X"F0",
		X"00",X"06",X"08",X"09",X"03",X"0D",X"08",X"06",X"02",X"04",X"01",X"08",X"02",X"06",X"05",X"04",
		X"09",X"09",X"09",X"0F",X"0F",X"00",X"0F",X"0F",X"0D",X"0D",X"0D",X"0D",X"0C",X"0E",X"07",X"03",
		X"00",X"00",X"08",X"08",X"09",X"09",X"09",X"09",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0B",X"0B",X"0B",X"0B",X"03",X"07",X"0E",X"0C",
		X"00",X"00",X"0F",X"0F",X"00",X"0E",X"0F",X"03",X"00",X"00",X"07",X"0F",X"0C",X"09",X"0B",X"0B",
		X"09",X"09",X"09",X"0F",X"0F",X"00",X"0F",X"0F",X"0D",X"0D",X"0D",X"0D",X"0C",X"0E",X"07",X"03",
		X"00",X"00",X"08",X"09",X"09",X"09",X"09",X"09",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"03",X"03",X"03",X"0F",X"0E",X"00",X"0F",X"0F",X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"0F",X"0F",
		X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"09",X"08",X"08",X"0F",X"0F",X"00",X"0F",X"0F",X"0D",X"0D",X"0D",X"0D",X"0C",X"0E",X"07",X"03",
		X"00",X"00",X"09",X"09",X"09",X"09",X"09",X"09",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"03",X"03",X"03",X"0F",X"0E",X"00",X"0F",X"0F",X"0B",X"00",X"00",X"0F",X"0F",X"00",X"0F",X"0F",
		X"00",X"00",X"0F",X"0F",X"00",X"0F",X"0F",X"03",X"00",X"00",X"0F",X"0F",X"08",X"0B",X"0B",X"0B",
		X"0C",X"0F",X"03",X"0C",X"07",X"01",X"00",X"00",X"0D",X"0E",X"07",X"01",X"00",X"00",X"00",X"00",
		X"01",X"0E",X"00",X"01",X"07",X"0C",X"03",X"0F",X"04",X"03",X"00",X"00",X"00",X"01",X"07",X"0E",
		X"03",X"00",X"00",X"0E",X"0F",X"01",X"0E",X"07",X"00",X"00",X"0F",X"07",X"08",X"0F",X"03",X"00",
		X"01",X"07",X"0C",X"03",X"0F",X"0F",X"03",X"03",X"00",X"00",X"03",X"0E",X"09",X"07",X"0E",X"00",
		X"00",X"00",X"80",X"C2",X"C2",X"C2",X"C0",X"C0",X"00",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"01",X"12",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"87",X"87",X"87",X"87",X"87",X"00",X"00",X"F0",X"F2",X"F3",X"71",X"70",X"30",X"00",X"00",
		X"F0",X"F0",X"F7",X"F6",X"F0",X"F0",X"03",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",
		X"00",X"00",X"87",X"87",X"87",X"87",X"87",X"C0",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",
		X"07",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C2",X"C2",X"C2",X"80",X"00",X"00",X"F2",X"F3",X"71",X"70",X"30",X"00",X"00",X"00",
		X"F0",X"F6",X"F7",X"F0",X"F0",X"10",X"03",X"06",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"00",
		X"00",X"00",X"80",X"C2",X"C2",X"CA",X"CC",X"CC",X"00",X"00",X"00",X"30",X"71",X"73",X"E2",X"E0",
		X"00",X"01",X"12",X"F0",X"FC",X"FC",X"56",X"16",X"0C",X"08",X"F0",X"F0",X"F3",X"F7",X"FF",X"FF",
		X"CC",X"8F",X"8F",X"8F",X"87",X"86",X"00",X"00",X"F0",X"F1",X"E2",X"62",X"71",X"30",X"00",X"00",
		X"96",X"9E",X"56",X"74",X"FC",X"F0",X"03",X"01",X"FF",X"FF",X"FF",X"F7",X"F3",X"F0",X"F0",X"0C",
		X"00",X"00",X"86",X"87",X"8F",X"8F",X"8F",X"CC",X"00",X"00",X"30",X"71",X"62",X"E2",X"F1",X"F0",
		X"07",X"01",X"F0",X"FC",X"74",X"56",X"9E",X"96",X"08",X"F0",X"F0",X"F3",X"F7",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CA",X"C2",X"C2",X"80",X"00",X"00",X"E0",X"E2",X"73",X"71",X"30",X"00",X"00",X"00",
		X"16",X"56",X"FC",X"FC",X"F0",X"10",X"03",X"06",X"FF",X"FF",X"F7",X"F3",X"F0",X"F0",X"08",X"00",
		X"0C",X"07",X"0B",X"81",X"48",X"0C",X"0E",X"C0",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"00",X"F0",X"C3",X"87",X"0F",X"F0",X"F0",X"01",X"E0",X"F0",X"1E",X"0F",X"0F",X"C3",X"F0",
		X"CC",X"CC",X"8C",X"8B",X"03",X"06",X"0C",X"00",X"70",X"71",X"31",X"30",X"10",X"00",X"00",X"00",
		X"FC",X"FE",X"32",X"32",X"F0",X"06",X"06",X"02",X"F3",X"F7",X"F7",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"08",X"81",X"83",X"87",X"83",X"00",X"00",X"30",X"70",X"70",X"E1",X"F0",X"F0",
		X"00",X"00",X"F0",X"C3",X"0F",X"0F",X"3C",X"F0",X"00",X"70",X"87",X"0F",X"0F",X"78",X"F0",X"F0",
		X"8B",X"8B",X"89",X"00",X"00",X"00",X"00",X"00",X"F1",X"F3",X"62",X"60",X"30",X"00",X"00",X"00",
		X"F8",X"FC",X"74",X"71",X"F1",X"0C",X"0C",X"08",X"F7",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"40",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"07",X"3C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"C0",X"C3",X"C3",X"C3",X"E1",X"F0",X"F0",
		X"00",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"F0",X"F4",X"F5",X"F1",X"F0",X"E1",X"40",X"00",
		X"F0",X"F0",X"F8",X"F8",X"F0",X"3C",X"07",X"00",X"F0",X"E1",X"C3",X"C3",X"C3",X"C0",X"08",X"00",
		X"00",X"80",X"C1",X"E1",X"E1",X"E1",X"E1",X"E0",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"30",
		X"0F",X"03",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"C1",X"80",X"00",X"00",X"30",X"31",X"11",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"FB",X"FB",X"F0",X"03",X"0F",X"00",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"08",X"00",
		X"00",X"00",X"82",X"CA",X"CE",X"CE",X"CC",X"CF",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"0F",X"12",X"F0",X"F7",X"CC",X"CC",X"E7",X"E1",X"08",X"F0",X"F0",X"F1",X"F3",X"7F",X"7F",X"7F",
		X"8F",X"8F",X"8F",X"8F",X"87",X"07",X"00",X"00",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",
		X"E7",X"CC",X"CC",X"F7",X"F0",X"12",X"0F",X"00",X"7F",X"7F",X"F3",X"F1",X"F0",X"F0",X"08",X"00",
		X"00",X"00",X"00",X"06",X"86",X"0E",X"8E",X"8E",X"00",X"00",X"00",X"30",X"71",X"73",X"F3",X"F1",
		X"00",X"01",X"07",X"F0",X"FC",X"30",X"12",X"9E",X"00",X"0E",X"E0",X"F0",X"F3",X"F7",X"FF",X"FF",
		X"88",X"88",X"8C",X"8C",X"84",X"04",X"00",X"00",X"F0",X"F1",X"F3",X"73",X"71",X"30",X"00",X"00",
		X"96",X"9E",X"12",X"30",X"FC",X"F0",X"07",X"01",X"FF",X"FF",X"FF",X"F7",X"F3",X"F0",X"E0",X"0E",
		X"08",X"0C",X"0F",X"0B",X"81",X"81",X"CC",X"CC",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"F0",
		X"00",X"30",X"30",X"70",X"F0",X"F0",X"E1",X"C3",X"01",X"C0",X"E0",X"E1",X"E1",X"F0",X"F0",X"79",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F3",X"F7",X"C4",X"40",X"30",X"01",X"01",
		X"C3",X"E9",X"E9",X"E9",X"EB",X"E3",X"09",X"03",X"79",X"3F",X"3F",X"2E",X"0C",X"0C",X"0C",X"08",
		X"00",X"08",X"0C",X"0F",X"83",X"81",X"85",X"8E",X"00",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"10",X"70",X"F0",X"F0",X"F0",X"C3",X"C3",X"40",X"E0",X"F0",X"E1",X"F0",X"F0",X"F0",X"79",
		X"8B",X"89",X"01",X"00",X"00",X"00",X"08",X"00",X"F3",X"F7",X"E6",X"62",X"30",X"01",X"01",X"00",
		X"E9",X"E9",X"61",X"71",X"F3",X"08",X"00",X"00",X"7B",X"3F",X"3F",X"0E",X"0E",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"F3",X"F7",X"C4",X"C0",X"E1",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"C0",X"C4",X"F7",X"F3",X"70",X"70",X"30",
		X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F4",X"F4",X"B0",X"B0",X"F4",X"B4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"F4",X"B0",X"B0",X"F4",X"F4",X"F0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F8",X"F8",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"F0",X"F0",X"F8",X"FD",X"F5",X"F1",X"F0",X"70",
		X"60",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F6",X"F6",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"70",X"F1",X"F3",X"F0",X"F0",X"70",X"30",X"00",
		X"F0",X"30",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"70",X"F3",X"F0",X"70",
		X"00",X"00",X"00",X"00",X"C3",X"BB",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"10",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"F2",X"F3",X"71",X"70",X"30",X"10",X"00",X"00",
		X"F0",X"F0",X"F7",X"F7",X"F0",X"F0",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F4",X"F6",X"F6",X"F2",X"70",X"30",X"00",X"F0",X"F0",X"F0",X"FE",X"FE",X"FC",X"F0",X"F0",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"10",X"30",X"71",X"71",X"F0",X"F0",
		X"00",X"70",X"F0",X"FE",X"FF",X"99",X"98",X"C3",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"F0",X"F0",X"71",X"71",X"30",X"10",X"00",X"00",
		X"C3",X"98",X"99",X"FF",X"FE",X"F0",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"30",X"71",X"F3",X"F3",X"E2",X"E0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"70",X"70",X"3C",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"E2",X"F3",X"F3",X"71",X"30",X"00",X"3C",X"70",X"70",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"F0",X"71",X"71",X"30",X"10",X"00",X"00",X"00",
		X"FE",X"FF",X"99",X"98",X"F0",X"16",X"02",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"F3",X"C0",X"C0",X"71",X"10",X"00",X"00",X"F8",X"FC",X"FC",X"FC",X"F8",X"F0",X"3C",X"08",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"30",X"70",X"F0",X"F4",X"FE",X"98",X"98",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"88",X"F0",X"F2",X"C4",X"C4",X"F7",X"F2",X"70",X"30",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"22",X"00",X"10",X"98",X"10",X"10",X"30",X"70",X"F2",X"F7",X"C4",X"C4",X"F2",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"98",X"10",X"00",X"00",X"22",X"00",X"00",X"98",X"98",X"FE",X"F4",X"F0",X"70",X"30",X"10",
		X"08",X"0C",X"06",X"C3",X"C3",X"F0",X"F0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"06",X"15",X"33",X"33",X"33",X"08",X"08",X"08",X"36",X"FE",X"FC",X"FC",X"F8",
		X"3C",X"3C",X"1E",X"1E",X"96",X"C3",X"E1",X"C1",X"00",X"00",X"22",X"01",X"88",X"88",X"11",X"11",
		X"33",X"30",X"3C",X"2C",X"20",X"30",X"10",X"00",X"F0",X"F0",X"FE",X"76",X"76",X"FC",X"F0",X"F0",
		X"0C",X"08",X"04",X"96",X"96",X"96",X"96",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"0F",X"0F",X"01",X"67",X"EF",X"FC",X"FC",X"F8",
		X"1E",X"1E",X"3C",X"78",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"89",X"88",X"00",X"00",X"44",X"44",
		X"33",X"30",X"3C",X"3D",X"31",X"B8",X"10",X"00",X"F0",X"F0",X"30",X"32",X"FE",X"FC",X"F0",X"F0",
		X"0E",X"C3",X"E9",X"ED",X"E5",X"E5",X"E1",X"E1",X"03",X"70",X"F3",X"F4",X"F4",X"F0",X"F0",X"F0",
		X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E1",X"E1",X"E1",X"E1",X"E5",X"E5",X"E8",X"C0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F6",X"F3",X"70",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F0",
		X"0E",X"CF",X"EF",X"EF",X"EF",X"EF",X"E7",X"E3",X"03",X"77",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"0F",X"FE",X"FC",X"F8",X"F0",X"0F",X"0F",X"0F",X"0F",X"FF",X"F7",X"F3",X"F1",X"1E",X"1E",X"1E",
		X"E1",X"E3",X"E7",X"EF",X"EF",X"EF",X"EE",X"CC",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"77",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"F8",X"FC",X"FE",X"1E",X"1E",X"1E",X"1E",X"F1",X"F3",X"F7",X"FF",
		X"00",X"00",X"81",X"0B",X"87",X"C1",X"C0",X"C0",X"00",X"07",X"00",X"30",X"70",X"F0",X"F0",X"F0",
		X"10",X"3C",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"84",X"83",X"03",X"01",X"01",X"00",X"00",X"00",X"F0",X"F4",X"F6",X"72",X"30",X"00",X"01",X"00",
		X"F0",X"F0",X"FC",X"FE",X"F0",X"03",X"0F",X"00",X"F0",X"F0",X"F0",X"C0",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"83",X"84",X"00",X"01",X"00",X"30",X"70",X"F0",X"F0",X"F0",
		X"00",X"0F",X"03",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"08",X"0C",X"C0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C1",X"87",X"0B",X"81",X"00",X"00",X"F0",X"F6",X"F2",X"70",X"30",X"00",X"07",X"00",
		X"F0",X"F0",X"F4",X"F6",X"F2",X"78",X"3C",X"10",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"88",X"77",X"00",X"77",X"88",X"88",X"EE",X"11",X"11",X"EE",X"00",X"EE",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"00",X"FF",X"44",X"00",X"00",X"00",X"EE",X"00",X"11",X"FF",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"88",X"77",X"00",X"77",X"88",X"88",X"EE",X"11",X"11",X"EE",X"00",X"EE",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"00",X"FF",X"44",X"22",X"11",X"00",X"EE",X"00",X"44",X"FF",X"44",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"77",X"00",X"77",X"88",X"77",X"00",X"EE",X"11",X"EE",X"00",X"EE",X"11",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"99",X"99",X"77",X"00",X"00",X"FF",X"44",X"EE",X"11",X"11",X"EE",X"00",X"11",X"FF",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"77",X"00",X"77",X"88",X"77",X"00",X"EE",X"11",X"EE",X"00",X"EE",X"11",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"88",X"44",X"66",X"99",X"99",X"44",X"11",X"99",X"55",X"33",X"EE",X"11",X"11",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"88",X"77",X"00",X"77",X"88",X"77",X"00",X"EE",X"11",X"EE",X"00",X"EE",X"11",X"EE",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"44",X"33",X"00",X"44",X"99",X"99",X"77",X"FF",X"44",X"44",X"CC",X"EE",X"11",X"11",X"EE",
		X"00",X"00",X"00",X"80",X"89",X"8B",X"8B",X"8B",X"00",X"00",X"30",X"73",X"E6",X"E2",X"F0",X"E6",
		X"00",X"00",X"F0",X"F8",X"35",X"3D",X"3D",X"35",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"83",X"81",X"80",X"0C",X"08",X"00",X"00",X"E6",X"F3",X"70",X"70",X"30",X"00",X"00",X"00",
		X"70",X"F8",X"0F",X"87",X"C3",X"30",X"00",X"00",X"EF",X"F0",X"F0",X"3C",X"0F",X"0F",X"00",X"00",
		X"08",X"88",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"30",
		X"01",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"3F",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"10",X"10",X"06",X"0F",X"3F",X"3F",X"0F",X"07",
		X"F0",X"F4",X"F6",X"F2",X"70",X"B8",X"FE",X"33",X"F0",X"F0",X"F0",X"FE",X"FE",X"FC",X"F0",X"F8",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"07",X"0F",X"3F",X"3F",X"0F",X"06",X"10",X"10",
		X"33",X"FE",X"B8",X"70",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"88",X"08",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"F4",X"F6",X"F2",X"F0",X"F0",X"70",X"30",X"01",X"F0",X"FE",X"FE",X"FC",X"F0",X"F0",X"F7",X"3F",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"30",X"70",X"71",X"F1",X"F0",X"F0",
		X"01",X"E1",X"F0",X"FE",X"FF",X"CC",X"CC",X"E1",X"0C",X"0E",X"E0",X"F0",X"F0",X"F0",X"F0",X"78",
		X"80",X"00",X"00",X"03",X"07",X"CF",X"07",X"00",X"F0",X"F1",X"F1",X"F0",X"70",X"30",X"00",X"00",
		X"EF",X"FF",X"CC",X"CC",X"F0",X"F0",X"F0",X"00",X"78",X"F0",X"F0",X"E0",X"E0",X"D1",X"FF",X"00",
		X"00",X"07",X"CF",X"07",X"03",X"80",X"80",X"C0",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"70",X"F0",X"F0",X"E6",X"EE",X"FF",X"F7",X"00",X"F7",X"D1",X"F0",X"70",X"70",X"F8",X"3C",
		X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",
		X"F0",X"E6",X"EE",X"FF",X"F7",X"F0",X"61",X"01",X"3C",X"70",X"70",X"F8",X"F0",X"F0",X"0E",X"0C",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"78",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"CC",X"F0",X"F0",X"F0",X"F0",X"F3",X"F7",X"F0",X"CB",
		X"2C",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C4",X"70",X"06",X"04",X"00",X"00",X"00",X"00",X"87",X"87",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"10",X"30",X"30",X"70",X"70",X"70",X"70",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"FE",X"32",X"30",X"F0",X"0C",X"09",X"03",X"03",X"FC",X"FC",X"FC",X"FC",X"CC",X"0E",X"0F",X"0F",
		X"00",X"80",X"00",X"40",X"C4",X"64",X"C0",X"20",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"E0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"00",X"F7",X"FF",X"FF",X"51",X"80",X"00",X"F0",X"F0",X"F2",X"F3",X"71",X"70",X"30",X"00",
		X"F0",X"F0",X"F0",X"F7",X"F6",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",
		X"00",X"80",X"51",X"FF",X"FF",X"F7",X"00",X"C0",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"20",X"C0",X"64",X"C4",X"40",X"00",X"80",X"00",X"F0",X"F2",X"F3",X"71",X"70",X"30",X"00",X"00",
		X"F0",X"F0",X"F7",X"F6",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"E0",X"00",
		X"00",X"80",X"40",X"B3",X"77",X"FF",X"77",X"F3",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"F7",X"CC",X"CC",X"F6",X"E1",X"00",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",X"78",
		X"20",X"C0",X"EC",X"C4",X"C0",X"CC",X"80",X"00",X"F0",X"F0",X"F1",X"F1",X"70",X"70",X"30",X"00",
		X"E1",X"98",X"98",X"FE",X"FC",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",X"F0",X"E0",X"F0",X"E0",X"F0",
		X"00",X"80",X"CC",X"C0",X"C4",X"EC",X"C0",X"20",X"00",X"30",X"70",X"70",X"F1",X"F1",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FC",X"FE",X"98",X"98",X"C3",X"F0",X"E0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"F3",X"77",X"FF",X"77",X"B3",X"40",X"80",X"00",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"00",X"00",
		X"C3",X"F4",X"CC",X"CC",X"F6",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"00",
		X"88",X"EE",X"33",X"91",X"51",X"A0",X"C0",X"A0",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"51",X"A0",X"D1",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"A0",X"C4",X"73",X"B3",X"66",X"CC",X"88",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",
		X"F0",X"F7",X"FF",X"99",X"90",X"F0",X"16",X"04",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"E0",X"11",
		X"00",X"00",X"80",X"40",X"80",X"51",X"F7",X"B3",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A0",X"D0",X"E0",X"F0",X"E0",X"F0",X"F0",X"F0",
		X"F3",X"B1",X"51",X"80",X"40",X"80",X"00",X"00",X"F0",X"F0",X"71",X"71",X"30",X"10",X"00",X"00",
		X"F0",X"FE",X"FF",X"32",X"30",X"F0",X"3C",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"00",X"00",X"70",X"F0",X"F3",X"F7",X"F7",X"F0",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F0",X"78",
		X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F7",X"F7",X"F3",X"F0",X"70",X"00",X"00",X"78",X"F0",X"F8",X"F8",X"F0",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"30",X"F0",X"F3",X"F7",X"F3",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F7",X"F3",X"F0",X"30",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"70",X"F3",X"F3",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F3",X"70",X"30",X"00",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"71",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"71",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"8F",X"0E",X"2E",X"3F",X"7F",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"00",
		X"89",X"01",X"30",X"62",X"E2",X"F1",X"F0",X"70",X"00",X"08",X"F1",X"75",X"74",X"E9",X"C3",X"87",
		X"F7",X"F7",X"F3",X"F3",X"F1",X"E0",X"00",X"0C",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"10",X"10",X"30",X"10",X"01",X"00",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"07",
		X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"77",X"77",X"FF",
		X"00",X"88",X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"77",X"33",X"33",X"33",X"11",
		X"00",X"01",X"01",X"30",X"71",X"62",X"E2",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F1",X"E2",X"62",X"71",X"30",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"0F",X"E1",X"F8",X"F8",X"BD",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"70",X"F3",X"C4",X"C4",X"F3",
		X"3D",X"3D",X"BD",X"F8",X"F8",X"E1",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"F3",X"C4",X"C4",X"F3",X"70",X"00",X"00",
		X"00",X"04",X"04",X"06",X"07",X"08",X"88",X"88",X"30",X"70",X"F3",X"F3",X"F1",X"F0",X"F0",X"F0",
		X"81",X"C3",X"21",X"30",X"FC",X"E1",X"C3",X"C3",X"00",X"01",X"03",X"8E",X"0E",X"3F",X"3F",X"7B",
		X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"70",X"70",X"30",X"10",X"00",X"00",X"00",X"00",
		X"C3",X"F0",X"F0",X"F0",X"F0",X"30",X"00",X"00",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"30",
		X"00",X"00",X"00",X"0E",X"03",X"CE",X"4E",X"6E",X"00",X"00",X"00",X"00",X"30",X"71",X"73",X"F1",
		X"00",X"00",X"00",X"00",X"F0",X"FC",X"21",X"03",X"00",X"00",X"00",X"02",X"0C",X"F3",X"F7",X"F7",
		X"6E",X"6E",X"EC",X"E0",X"E0",X"E0",X"C0",X"80",X"F0",X"F3",X"F3",X"F1",X"70",X"70",X"10",X"00",
		X"C3",X"21",X"30",X"FC",X"E1",X"E1",X"F0",X"00",X"E7",X"C3",X"87",X"0F",X"1E",X"3C",X"F0",X"F0",
		X"01",X"0F",X"0B",X"81",X"C8",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"0F",X"01",X"01",X"F0",X"90",X"98",X"EF",X"E1",X"08",X"08",X"78",X"F0",X"F1",X"7B",X"7B",X"7B",
		X"CC",X"CC",X"CC",X"C8",X"81",X"0B",X"0F",X"01",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"E7",X"98",X"98",X"F6",X"F0",X"01",X"01",X"0F",X"7B",X"7B",X"F3",X"F1",X"F0",X"78",X"08",X"08",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"01",X"00",X"00",X"00",X"00",X"30",X"71",X"73",X"F3",X"F1",
		X"07",X"06",X"16",X"F0",X"FC",X"30",X"12",X"9E",X"0E",X"00",X"E0",X"F0",X"F6",X"FF",X"FF",X"FF",
		X"00",X"01",X"0F",X"03",X"01",X"00",X"00",X"00",X"F0",X"F3",X"F3",X"71",X"30",X"00",X"00",X"00",
		X"96",X"9E",X"12",X"30",X"F0",X"16",X"06",X"07",X"FF",X"FF",X"FF",X"F6",X"F0",X"E0",X"00",X"0E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"FF",X"7F",X"0F",X"0F",X"0F",X"87",X"C3",X"E1",X"F7",X"C3",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F3",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F3",X"F7",
		X"97",X"87",X"C3",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"F0",X"F1",X"F1",X"F3",X"F3",X"E1",X"E1",X"F0",
		X"F0",X"F0",X"F0",X"F1",X"F1",X"F3",X"F7",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"4F",X"4F",X"4F",X"4F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"2F",X"0F",X"8F",X"FF",X"9F",X"8F",X"CF",X"CF",X"CF",X"DF",X"5F",
		X"5F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",X"5F",X"5F",X"5F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"2F",X"0F",X"0F",X"B5",X"A5",X"A5",X"A5",X"87",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"E7",X"F7",X"B7",X"B7",X"B5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F1",X"F1",X"F3",X"F3",X"F7",X"F7",X"F7",
		X"F1",X"F1",X"F1",X"F3",X"F3",X"F7",X"F7",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F1",X"F3",X"C3",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"B7",X"B7",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"0F",X"0F",X"87",X"C3",X"E1",X"E1",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"0F",X"FF",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"8F",X"CF",X"CF",X"EF",X"FF",X"FF",X"E1",X"F3",X"F3",X"F3",X"F7",X"F7",X"FF",X"FF",
		X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"2F",X"0F",X"0F",X"87",X"87",X"C3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F3",
		X"F1",X"F1",X"F3",X"F3",X"F7",X"F7",X"F7",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C3",X"C3",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F7",X"FF",X"FF",X"FF",X"1F",X"0F",X"87",X"87",X"F0",X"F0",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F1",X"F1",X"F3",X"F3",X"F3",X"F7",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"B4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"87",X"87",X"C3",X"C3",X"E1",X"F0",X"F0",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",
		X"8F",X"8F",X"EF",X"AF",X"1F",X"0F",X"0F",X"0F",X"3F",X"1F",X"1F",X"0F",X"87",X"87",X"87",X"A5",
		X"7F",X"7F",X"1F",X"8F",X"CF",X"EF",X"FF",X"FF",X"AF",X"CF",X"EF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"1F",X"1F",X"9F",X"DF",X"FF",X"FF",X"FF",X"FF",X"8F",X"8F",X"CF",X"CF",X"EF",X"FF",X"FF",X"6F",
		X"FF",X"9F",X"1F",X"9F",X"DF",X"5F",X"3F",X"3F",X"3F",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"8F",X"8F",X"0F",
		X"CF",X"EF",X"EF",X"7F",X"7F",X"3F",X"1F",X"FF",X"DF",X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"9F",X"8F",X"87",X"C7",X"E7",X"E7",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F3",X"F3",X"F3",X"F7",X"F7",X"F7",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"9F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"AF",X"EF",X"EF",X"6F",X"6F",X"2F",X"8F",X"8F",X"9F",X"8F",X"CF",X"CF",X"EF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"EF",X"EF",X"6F",X"6F",X"2F",X"2F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2F",
		X"FF",X"FF",X"7F",X"BF",X"9F",X"4F",X"0F",X"0F",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"2F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"3F",X"7F",X"7F",X"FF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",
		X"FF",X"BF",X"BF",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D3",X"F1",X"F3",X"F3",X"F7",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",
		X"7F",X"3F",X"BF",X"BF",X"BF",X"BF",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"1F",X"1F",X"8F",X"8F",X"CF",X"EF",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"5F",X"7F",X"3F",X"1F",X"1F",X"0F",X"1F",
		X"3F",X"BF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"9F",X"CF",X"6F",X"6F",X"3F",X"BF",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"9F",X"FF",X"7F",X"FF",X"FF",X"FF",X"3F",X"0F",X"1F",X"0F",X"8F",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"CF",X"8F",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"CF",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"0F",X"0F",X"0F",X"0F",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",
		X"8F",X"8F",X"9F",X"9F",X"9F",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"CF",X"CF",X"8F",X"8F",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"DF",X"DF",X"DF",X"CF",X"CF",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"8F",X"9F",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"2F",X"2F",X"2F",X"2F",X"0F",X"0F",X"0F",X"0F",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"6F",X"6F",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"8F",X"8F",X"AF",X"AF",X"AF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"DF",X"CF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"3F",X"3F",X"1F",X"9F",X"9F",X"9F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"3F",X"CF",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"1F",X"1F",X"1F",X"1F",X"8F",X"8F",X"8F",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"BF",X"BF",X"BF",X"9F",X"DF",X"DF",X"DF",X"DF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"2F",X"2F",X"2F",X"2F",X"3F",X"3F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"9F",X"FF",X"9F",X"DF",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"CF",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"3D",X"3D",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"1E",X"1E",X"1E",X"1E",X"3C",X"3C",X"3D",X"3D",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"3D",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"EF",X"CF",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"CF",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"CF",X"CF",X"CF",X"CF",
		X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"1E",X"1E",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"CF",X"EF",X"EF",X"EF",
		X"F7",X"F7",X"F3",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F3",X"F3",X"F1",X"F1",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"8F",X"CF",X"CF",X"EF",X"EF",X"0F",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"3C",X"1E",X"1E",X"0F",X"3C",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"78",X"78",X"3C",X"3C",
		X"F7",X"F7",X"F7",X"F7",X"F3",X"F3",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"F3",X"F3",X"F3",X"F3",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"EF",X"0F",X"8F",X"8F",X"CF",X"CF",X"EF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"3C",X"3C",X"78",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F3",X"F1",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"EF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"CF",X"CF",X"EF",X"EF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"3C",X"F0",X"F0",X"78",X"78",X"3C",X"1E",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"1E",X"1E",X"1E",X"3C",X"78",X"8F",X"8F",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"CF",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",
		X"8F",X"8F",X"8F",X"9F",X"9F",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CF",X"CF",X"CF",X"EF",X"EF",X"EF",X"FF",X"FF",
		X"78",X"78",X"3C",X"3C",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",X"8F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"3C",X"3C",X"1E",X"1E",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"3C",X"3C",X"3C",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",
		X"3C",X"3C",X"3C",X"3C",X"78",X"78",X"78",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"78",X"78",X"78",X"78",X"3C",X"3C",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",
		X"F0",X"C7",X"C7",X"E7",X"EF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"78",X"78",X"79",X"79",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"9F",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F1",X"F1",X"F3",X"F3",X"F3",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"F3",X"F7",X"F7",X"F7",X"FF",X"FF",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F3",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F3",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"8F",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"8F",X"8F",X"8F",X"8F",X"8F",X"CF",X"CF",X"CF",
		X"F3",X"F3",X"F3",X"7B",X"3F",X"7F",X"7F",X"7F",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",
		X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F3",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"3C",X"3C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"F3",X"F3",X"F7",X"F7",X"F7",X"F7",
		X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F1",
		X"F1",X"F1",X"F3",X"F3",X"F3",X"F7",X"F7",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F3",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F3",
		X"FF",X"FF",X"FF",X"F7",X"F3",X"F3",X"F1",X"F1",X"F7",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"F7",X"F3",X"F3",X"F7",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"4F",X"0F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",
		X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"B4",X"F0",X"F0",X"B4",X"B4",X"A5",X"A5",X"A5",X"A5",
		X"0F",X"2D",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"2D",X"A5",X"A5",X"A5",X"A5",
		X"5F",X"5F",X"5F",X"5F",X"4F",X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"0F",X"0F",
		X"FF",X"DF",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"DF",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"7F",X"FF",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"A5",X"A5",X"2D",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",X"5F",X"5F",X"5F",X"7F",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",X"5F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",
		X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"B4",X"A5",X"A5",X"A5",X"A5",X"F0",X"B4",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"B4",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"B4",
		X"5F",X"4F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",X"5F",X"5F",X"4F",X"4F",X"0F",
		X"5F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"1F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"0F",X"0F",X"0F",X"1F",X"5F",X"5F",X"5F",X"5F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"A5",X"A5",
		X"A5",X"B4",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"B4",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"2D",X"2D",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",X"2D",
		X"FF",X"FF",X"DF",X"DF",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"7F",X"FF",X"FF",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"7F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"5F",X"5F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",
		X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",X"F0",X"B4",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"A5",X"B4",X"B4",X"F0",X"F0",X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",X"B4",X"B4",X"F0",
		X"2D",X"2D",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",X"2D",X"2D",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2D",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",X"5F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"2D",X"2D",X"2D",X"A5",X"A5",X"A5",X"A5",
		X"0F",X"0F",X"0F",X"2D",X"2D",X"2D",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"5F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"7F",X"7F",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A5",X"A5",X"B4",X"B4",X"B4",X"B4",X"F0",X"F0",
		X"B4",X"B4",X"B4",X"B4",X"B4",X"B4",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"2D",X"2D",X"2D",X"2D",
		X"0F",X"0F",X"0F",X"0F",X"2D",X"2D",X"2D",X"2D",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"5F",X"5F",X"4F",X"4F",X"4F",X"4F",X"0F",X"0F",
		X"5F",X"5F",X"4F",X"4F",X"4F",X"4F",X"0F",X"0F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",
		X"DF",X"DF",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"E1",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"F0",X"F0",X"E1",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"B4",X"B4",X"B4",X"B4",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"B4",X"B4",X"B4",X"B4",
		X"B4",X"B4",X"B4",X"B4",X"F0",X"F0",X"F0",X"F0",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"A5",X"A5",X"A5",X"A5",X"B4",X"B4",X"B4",X"B4",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"5F",X"5F",X"4F",X"4F",X"4F",X"4F",X"0F",X"0F",X"FF",X"DF",X"DF",X"DF",X"5F",X"5F",X"5F",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"DF",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"A5",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"87",X"E1",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"A5",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"A5",X"A5",X"A5",X"A5",X"B4",X"B4",X"B4",X"B4",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"A5",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"5F",X"5F",X"5F",X"5F",X"5F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"5F",
		X"CF",X"CF",X"CF",X"CF",X"8F",X"8F",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"C2",X"C2",X"C2",X"C0",X"C0",X"00",X"00",X"00",X"30",X"60",X"40",X"D1",X"F1",
		X"00",X"01",X"12",X"F0",X"30",X"30",X"9A",X"9E",X"0C",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"87",X"87",X"87",X"87",X"86",X"00",X"00",X"F0",X"E0",X"D1",X"51",X"60",X"30",X"00",X"00",
		X"96",X"16",X"9A",X"B8",X"30",X"F0",X"03",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",
		X"00",X"00",X"86",X"87",X"87",X"87",X"87",X"C0",X"00",X"00",X"30",X"60",X"51",X"D1",X"E0",X"F0",
		X"07",X"01",X"F0",X"30",X"B8",X"9A",X"16",X"96",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C2",X"C2",X"C2",X"80",X"00",X"00",X"F1",X"D1",X"40",X"60",X"30",X"00",X"00",X"00",
		X"9E",X"9A",X"30",X"30",X"F0",X"10",X"03",X"06",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"00",
		X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"80",X"00",X"00",X"00",X"10",X"30",X"20",X"60",X"70",
		X"00",X"00",X"01",X"F0",X"30",X"10",X"DC",X"DE",X"00",X"0C",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"0E",X"0E",X"0E",X"0C",X"00",X"00",X"00",X"70",X"70",X"60",X"20",X"30",X"10",X"00",X"00",
		X"96",X"16",X"DE",X"DC",X"30",X"F0",X"01",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"0C",
		X"00",X"00",X"00",X"0C",X"0E",X"0E",X"0E",X"80",X"00",X"00",X"10",X"30",X"20",X"60",X"70",X"70",
		X"07",X"01",X"F0",X"30",X"DC",X"DE",X"16",X"96",X"00",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"84",X"84",X"84",X"00",X"00",X"00",X"00",X"70",X"60",X"20",X"30",X"10",X"00",X"00",X"00",
		X"DE",X"DC",X"10",X"30",X"F0",X"03",X"06",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"00",X"00",X"01",X"12",X"F0",X"90",X"76",X"45",X"00",X"00",X"0C",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"C3",X"45",X"76",X"90",X"F0",X"12",X"01",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"80",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"00",X"07",X"12",X"F0",X"90",X"76",X"45",X"C3",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"84",X"84",X"84",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"45",X"76",X"90",X"F0",X"12",X"07",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"01",X"F0",X"90",X"A3",X"00",X"00",X"00",X"08",X"00",X"F0",X"F0",X"F0",
		X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"A3",X"90",X"F0",X"01",X"00",X"00",X"00",X"F0",X"E1",X"E1",X"E1",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"02",X"01",X"F0",X"90",X"A3",X"E1",X"00",X"00",X"00",X"00",X"E1",X"E1",X"E1",X"F0",
		X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A3",X"90",X"F0",X"01",X"02",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"70",X"F0",X"00",X"00",X"00",X"00",X"08",X"00",X"E1",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"A0",X"70",X"01",X"00",X"00",X"00",X"00",X"E0",X"C3",X"C3",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"01",X"70",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"C3",X"C3",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"70",X"01",X"02",X"00",X"00",X"00",X"00",X"E1",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"C2",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"30",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"30",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C2",X"C2",X"C2",X"C0",X"C0",X"00",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"01",X"12",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"87",X"87",X"87",X"87",X"87",X"00",X"00",X"F0",X"D0",X"C0",X"60",X"70",X"30",X"00",X"00",
		X"F0",X"F0",X"80",X"90",X"F0",X"F0",X"03",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",
		X"00",X"00",X"87",X"87",X"87",X"87",X"87",X"C0",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",
		X"07",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C2",X"C2",X"C2",X"80",X"00",X"00",X"D0",X"C0",X"60",X"70",X"30",X"00",X"00",X"00",
		X"F0",X"90",X"80",X"F0",X"F0",X"10",X"03",X"06",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"00",
		X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"00",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"0C",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"70",X"60",X"60",X"30",X"30",X"10",X"00",X"00",
		X"F0",X"F0",X"40",X"40",X"F0",X"F0",X"01",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"0C",
		X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"80",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"07",X"01",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"84",X"84",X"84",X"00",X"00",X"00",X"00",X"60",X"60",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F0",X"40",X"40",X"F0",X"F0",X"03",X"06",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"84",X"84",X"84",X"80",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"00",X"00",X"01",X"12",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"0C",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"70",X"40",X"C0",X"F0",X"F0",X"12",X"01",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"80",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"00",X"07",X"12",X"F0",X"F0",X"F0",X"F0",X"70",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"84",X"84",X"84",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"F0",X"F0",X"12",X"07",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"01",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"08",X"00",X"F0",X"F0",X"F0",
		X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"50",X"C0",X"F0",X"01",X"00",X"00",X"00",X"F0",X"E1",X"E1",X"E1",X"00",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"02",X"01",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"E1",X"E1",X"E1",X"F0",
		X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"C0",X"F0",X"01",X"02",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"07",X"0B",X"81",X"48",X"0C",X"0E",X"C0",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"00",X"F0",X"C3",X"87",X"0F",X"F0",X"F0",X"01",X"E0",X"F0",X"1E",X"0F",X"0F",X"C3",X"F0",
		X"C0",X"C0",X"84",X"83",X"03",X"06",X"0C",X"00",X"70",X"60",X"20",X"30",X"10",X"00",X"00",X"00",
		X"30",X"10",X"DC",X"DC",X"F0",X"06",X"06",X"02",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"08",X"81",X"83",X"87",X"83",X"00",X"00",X"30",X"70",X"70",X"E1",X"F0",X"F0",
		X"00",X"00",X"F0",X"C3",X"0F",X"0F",X"3C",X"F0",X"00",X"70",X"87",X"0F",X"0F",X"78",X"F0",X"F0",
		X"83",X"83",X"81",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"51",X"71",X"30",X"00",X"00",X"00",
		X"70",X"30",X"B8",X"B8",X"F0",X"0C",X"0C",X"08",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"08",X"06",X"0A",X"80",X"08",X"0C",X"80",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"00",X"00",X"00",X"F0",X"C3",X"87",X"F0",X"F0",X"00",X"01",X"E0",X"F0",X"1E",X"0F",X"87",X"F0",
		X"80",X"80",X"08",X"06",X"0C",X"08",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"90",X"76",X"76",X"F0",X"06",X"02",X"00",X"00",X"F0",X"F0",X"F0",X"E0",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"08",X"02",X"06",X"0E",X"06",X"00",X"00",X"00",X"10",X"30",X"70",X"70",X"70",
		X"00",X"00",X"00",X"F0",X"C3",X"0F",X"1E",X"F0",X"00",X"00",X"E0",X"0F",X"0F",X"3C",X"F0",X"F0",
		X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"60",X"20",X"10",X"00",X"00",X"00",X"00",
		X"30",X"FC",X"FC",X"F0",X"0C",X"08",X"00",X"00",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"04",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"F0",X"C3",X"87",X"F0",X"00",X"00",X"03",X"C0",X"E1",X"1E",X"0F",X"F0",
		X"00",X"00",X"0C",X"0C",X"08",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"D4",X"F0",X"06",X"02",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"F0",X"87",X"0F",X"F0",X"00",X"00",X"00",X"C0",X"0F",X"2C",X"E0",X"E1",
		X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"30",X"B8",X"F0",X"0C",X"08",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"E1",X"C3",X"F0",X"00",X"00",X"00",X"C3",X"E1",X"1E",X"0F",X"F0",
		X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E2",X"70",X"02",X"01",X"00",X"00",X"00",X"F0",X"F0",X"E1",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"F0",X"C3",X"87",X"F0",X"00",X"00",X"00",X"C0",X"0E",X"2C",X"E0",X"E1",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"D4",X"F0",X"04",X"04",X"00",X"00",X"00",X"E1",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"10",X"30",X"60",X"60",X"F0",X"F0",
		X"00",X"70",X"F0",X"10",X"00",X"66",X"76",X"C3",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"F0",X"F0",X"60",X"60",X"30",X"10",X"00",X"00",
		X"C3",X"76",X"66",X"00",X"10",X"F0",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"30",X"60",X"C0",X"C0",X"D1",X"D1",X"F0",X"F0",X"F0",X"70",X"70",X"70",X"F8",X"F8",X"3C",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"D1",X"D1",X"C0",X"C0",X"60",X"30",X"00",X"3C",X"F8",X"F8",X"70",X"70",X"70",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"10",X"30",X"20",X"70",X"70",
		X"00",X"00",X"70",X"F0",X"10",X"66",X"76",X"C3",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"20",X"30",X"10",X"00",X"00",X"00",
		X"C3",X"76",X"66",X"10",X"F0",X"70",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"60",X"40",X"D1",X"D1",X"F0",X"00",X"F0",X"F0",X"70",X"70",X"F8",X"F8",X"3C",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"D1",X"D1",X"40",X"60",X"30",X"00",X"00",X"3C",X"F8",X"F8",X"70",X"70",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",
		X"00",X"00",X"00",X"70",X"90",X"76",X"54",X"C3",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"C3",X"54",X"76",X"90",X"70",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"20",X"51",X"51",X"70",X"00",X"00",X"F0",X"F0",X"70",X"F8",X"70",X"3C",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"51",X"51",X"20",X"30",X"00",X"00",X"00",X"3C",X"70",X"F8",X"70",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"70",X"B0",X"54",X"D2",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D2",X"54",X"B0",X"70",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"20",X"20",X"30",X"00",X"00",X"00",X"F0",X"F0",X"70",X"F8",X"B4",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"B4",X"F8",X"70",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"D0",X"70",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"70",X"70",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"10",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"D0",X"C0",X"60",X"70",X"30",X"10",X"00",X"00",
		X"F0",X"F0",X"80",X"80",X"F0",X"F0",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"B0",X"90",X"90",X"D0",X"70",X"30",X"00",X"F0",X"F0",X"F0",X"10",X"10",X"30",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F0",X"40",X"40",X"F0",X"F0",X"70",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"D0",X"C0",X"40",X"60",X"30",X"00",X"00",X"F0",X"F0",X"90",X"90",X"90",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",
		X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"70",X"40",X"D0",X"F0",X"70",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"30",X"70",X"70",X"70",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"60",X"60",X"30",X"30",X"00",X"00",X"00",X"F0",X"F0",X"90",X"90",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"C0",X"F0",X"70",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"20",X"30",X"10",X"00",X"00",X"00",X"00",X"F0",X"B0",X"90",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",
		X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"F0",X"60",X"60",X"30",X"10",X"00",X"00",X"00",
		X"10",X"00",X"66",X"76",X"F0",X"16",X"02",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"F3",X"F3",X"60",X"10",X"00",X"00",X"70",X"30",X"30",X"30",X"70",X"F0",X"3C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"00",X"70",X"F0",X"F0",X"F0",X"F0",X"90",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"66",X"F6",X"F0",X"16",X"02",X"00",X"00",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"70",X"70",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"71",X"71",X"30",X"10",X"00",X"00",X"00",X"30",X"B8",X"B8",X"70",X"F0",X"3C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",
		X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"90",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"D4",X"F0",X"16",X"02",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"30",X"B8",X"B8",X"F0",X"3C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"30",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"F0",X"34",X"04",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"30",X"B8",X"F0",X"78",X"08",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
